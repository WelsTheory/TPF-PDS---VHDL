library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sin_entity is
    Port (
        address: in std_logic_vector(11 downto 0);
        sine: out std_logic_vector(15 downto 0)
    );
end entity;

architecture Behavioral of sin_entity is
    
    type mem is array(0 to 4095) of real;
    constant my_rom: mem := (
0=>750.0,
1=>751.1507660882452,
2=>752.3015294673039,
3=>753.4522874279961,
4=>754.6030372611546,
5=>755.753776257631,
6=>756.9045017083026,
7=>758.0552109040789,
8=>759.2059011359072,
9=>760.3565696947796,
10=>761.5072138717394,
11=>762.657830957887,
12=>763.8084182443869,
13=>764.9589730224735,
14=>766.1094925834578,
15=>767.2599742187339,
16=>768.4104152197849,
17=>769.5608128781896,
18=>770.7111644856291,
19=>771.8614673338926,
20=>773.0117187148844,
21=>774.1619159206297,
22=>775.3120562432812,
23=>776.4621369751259,
24=>777.6121554085908,
25=>778.7621088362494,
26=>779.9119945508287,
27=>781.0618098452147,
28=>782.2115520124596,
29=>783.3612183457872,
30=>784.5108061386004,
31=>785.6603126844866,
32=>786.8097352772246,
33=>787.9590712107911,
34=>789.1083177793663,
35=>790.2574722773412,
36=>791.4065319993234,
37=>792.5554942401438,
38=>793.7043562948625,
39=>794.8531154587756,
40=>796.0017690274216,
41=>797.1503142965872,
42=>798.2987485623146,
43=>799.4470691209068,
44=>800.5952732689349,
45=>801.7433583032437,
46=>802.8913215209587,
47=>804.0391602194923,
48=>805.1868716965495,
49=>806.3344532501353,
50=>807.4819021785605,
51=>808.629215780448,
52=>809.7763913547393,
53=>810.9234262007011,
54=>812.070317617931,
55=>813.2170629063646,
56=>814.3636593662814,
57=>815.5101042983111,
58=>816.6563950034406,
59=>817.8025287830194,
60=>818.9485029387668,
61=>820.0943147727776,
62=>821.2399615875289,
63=>822.3854406858864,
64=>823.5307493711103,
65=>824.6758849468624,
66=>825.8208447172119,
67=>826.9656259866418,
68=>828.1102260600554,
69=>829.2546422427824,
70=>830.3988718405859,
71=>831.5429121596676,
72=>832.6867605066755,
73=>833.830414188709,
74=>834.973870513326,
75=>836.1171267885493,
76=>837.260180322872,
77=>838.4030284252652,
78=>839.5456684051833,
79=>840.6880975725705,
80=>841.8303132378678,
81=>842.9723127120184,
82=>844.1140933064745,
83=>845.255652333204,
84=>846.396987104696,
85=>847.5380949339676,
86=>848.6789731345704,
87=>849.8196190205964,
88=>850.9600299066846,
89=>852.1002031080272,
90=>853.2401359403761,
91=>854.3798257200491,
92=>855.5192697639359,
93=>856.658465389505,
94=>857.7974099148097,
95=>858.9361006584944,
96=>860.074534939801,
97=>861.212710078575,
98=>862.3506233952725,
99=>863.4882722109653,
100=>864.6256538473483,
101=>865.7627656267455,
102=>866.8996048721159,
103=>868.0361689070603,
104=>869.1724550558274,
105=>870.3084606433201,
106=>871.4441829951019,
107=>872.5796194374028,
108=>873.7147672971263,
109=>874.8496239018549,
110=>875.9841865798571,
111=>877.1184526600933,
112=>878.2524194722221,
113=>879.3860843466066,
114=>880.519444614321,
115=>881.6524976071563,
116=>882.785240657627,
117=>883.9176710989775,
118=>885.0497862651878,
119=>886.1815834909803,
120=>887.313060111826,
121=>888.4442134639506,
122=>889.5750408843409,
123=>890.7055397107508,
124=>891.8357072817082,
125=>892.9655409365205,
126=>894.0950380152813,
127=>895.2241958588768,
128=>896.3530118089915,
129=>897.481483208115,
130=>898.6096073995482,
131=>899.737381727409,
132=>900.8648035366396,
133=>901.9918701730112,
134=>903.1185789831321,
135=>904.2449273144524,
136=>905.3709125152711,
137=>906.4965319347423,
138=>907.6217829228806,
139=>908.7466628305685,
140=>909.8711690095621,
141=>910.9952988124971,
142=>912.1190495928956,
143=>913.2424187051718,
144=>914.3654035046382,
145=>915.4880013475126,
146=>916.6102095909235,
147=>917.7320255929166,
148=>918.853446712461,
149=>919.9744703094558,
150=>921.0950937447354,
151=>922.2153143800767,
152=>923.3351295782047,
153=>924.454536702799,
154=>925.5735331184999,
155=>926.6921161909145,
156=>927.8102832866232,
157=>928.9280317731855,
158=>930.0453590191464,
159=>931.162262394043,
160=>932.2787392684097,
161=>933.3947870137856,
162=>934.5104030027196,
163=>935.6255846087772,
164=>936.7403292065467,
165=>937.854634171645,
166=>938.9684968807242,
167=>940.0819147114772,
168=>941.194885042645,
169=>942.3074052540212,
170=>943.41947272646,
171=>944.5310848418807,
172=>945.6422389832749,
173=>946.7529325347126,
174=>947.863162881348,
175=>948.9729274094256,
176=>950.0822235062867,
177=>951.1910485603755,
178=>952.2993999612451,
179=>953.4072750995635,
180=>954.5146713671203,
181=>955.6215861568322,
182=>956.7280168627494,
183=>957.8339608800619,
184=>958.9394156051055,
185=>960.0443784353679,
186=>961.1488467694944,
187=>962.2528180072954,
188=>963.3562895497507,
189=>964.459258799017,
190=>965.5617231584331,
191=>966.663680032527,
192=>967.7651268270212,
193=>968.8660609488387,
194=>969.9664798061099,
195=>971.0663808081781,
196=>972.1657613656059,
197=>973.2646188901809,
198=>974.3629507949222,
199=>975.4607544940864,
200=>976.5580274031734,
201=>977.6547669389329,
202=>978.7509705193702,
203=>979.8466355637527,
204=>980.941759492615,
205=>982.0363397277662,
206=>983.130373692295,
207=>984.2238588105765,
208=>985.3167925082778,
209=>986.4091722123638,
210=>987.5009953511044,
211=>988.5922593540789,
212=>989.6829616521838,
213=>990.7730996776372,
214=>991.8626708639864,
215=>992.9516726461127,
216=>994.0401024602377,
217=>995.1279577439303,
218=>996.2152359361114,
219=>997.3019344770605,
220=>998.3880508084223,
221=>999.4735823732115,
222=>1000.5585266158198,
223=>1001.6428809820216,
224=>1002.72664291898,
225=>1003.8098098752529,
226=>1004.8923793007986,
227=>1005.9743486469824,
228=>1007.0557153665826,
229=>1008.1364769137957,
230=>1009.2166307442432,
231=>1010.2961743149772,
232=>1011.3751050844867,
233=>1012.4534205127032,
234=>1013.531118061007,
235=>1014.6081951922329,
236=>1015.6846493706764,
237=>1016.7604780620995,
238=>1017.835678733737,
239=>1018.9102488543019,
240=>1019.9841858939917,
241=>1021.0574873244947,
242=>1022.130150618995,
243=>1023.2021732521796,
244=>1024.2735527002433,
245=>1025.3442864408958,
246=>1026.4143719533658,
247=>1027.4838067184091,
248=>1028.5525882183133,
249=>1029.6207139369037,
250=>1030.6881813595496,
251=>1031.7549879731703,
252=>1032.8211312662404,
253=>1033.8866087287963,
254=>1034.951417852442,
255=>1036.015556130355,
256=>1037.079021057292,
257=>1038.141810129595,
258=>1039.203920845197,
259=>1040.265350703628,
260=>1041.3260972060211,
261=>1042.3861578551182,
262=>1043.4455301552755,
263=>1044.5042116124705,
264=>1045.562199734306,
265=>1046.6194920300184,
266=>1047.676086010481,
267=>1048.7319791882119,
268=>1049.7871690773786,
269=>1050.841653193805,
270=>1051.8954290549757,
271=>1052.948494180043,
272=>1054.000846089833,
273=>1055.0524823068502,
274=>1056.103400355284,
275=>1057.1535977610154,
276=>1058.2030720516207,
277=>1059.2518207563796,
278=>1060.29984140628,
279=>1061.3471315340228,
280=>1062.3936886740298,
281=>1063.4395103624481,
282=>1064.484594137156,
283=>1065.5289375377693,
284=>1066.5725381056468,
285=>1067.615393383896,
286=>1068.657500917379,
287=>1069.698858252718,
288=>1070.7394629383025,
289=>1071.7793125242924,
290=>1072.8184045626263,
291=>1073.8567366070256,
292=>1074.8943062130015,
293=>1075.93111093786,
294=>1076.9671483407076,
295=>1078.0024159824575,
296=>1079.0369114258347,
297=>1080.070632235383,
298=>1081.1035759774688,
299=>1082.1357402202887,
300=>1083.1671225338741,
301=>1084.1977204900973,
302=>1085.2275316626774,
303=>1086.2565536271852,
304=>1087.2847839610502,
305=>1088.312220243565,
306=>1089.3388600558922,
307=>1090.3647009810686,
308=>1091.389740604013,
309=>1092.4139765115294,
310=>1093.4374062923148,
311=>1094.4600275369637,
312=>1095.4818378379741,
313=>1096.5028347897533,
314=>1097.5230159886232,
315=>1098.5423790328264,
316=>1099.5609215225313,
317=>1100.5786410598387,
318=>1101.5955352487863,
319=>1102.611601695355,
320=>1103.6268380074744,
321=>1104.6412417950282,
322=>1105.654810669861,
323=>1106.667542245782,
324=>1107.679434138572,
325=>1108.6904839659887,
326=>1109.7006893477717,
327=>1110.7100479056494,
328=>1111.7185572633432,
329=>1112.7262150465742,
330=>1113.733018883068,
331=>1114.738966402561,
332=>1115.7440552368046,
333=>1116.7482830195731,
334=>1117.751647386667,
335=>1118.7541459759198,
336=>1119.755776427203,
337=>1120.7565363824326,
338=>1121.7564234855731,
339=>1122.7554353826445,
340=>1123.753569721727,
341=>1124.7508241529667,
342=>1125.7471963285816,
343=>1126.7426839028662,
344=>1127.7372845321984,
345=>1128.730995875043,
346=>1129.7238155919592,
347=>1130.7157413456055,
348=>1131.7067708007444,
349=>1132.6969016242488,
350=>1133.6861314851076,
351=>1134.6744580544296,
352=>1135.6618790054515,
353=>1136.6483920135413,
354=>1137.6339947562046,
355=>1138.6186849130906,
356=>1139.6024601659958,
357=>1140.5853181988716,
358=>1141.5672566978285,
359=>1142.5482733511412,
360=>1143.528365849256,
361=>1144.5075318847935,
362=>1145.485769152556,
363=>1146.4630753495326,
364=>1147.4394481749036,
365=>1148.414885330048,
366=>1149.389384518546,
367=>1150.3629434461873,
368=>1151.3355598209744,
369=>1152.3072313531293,
370=>1153.2779557550982,
371=>1154.2477307415568,
372=>1155.2165540294166,
373=>1156.184423337829,
374=>1157.1513363881916,
375=>1158.1172909041534,
376=>1159.0822846116196,
377=>1160.0463152387576,
378=>1161.0093805160025,
379=>1161.9714781760615,
380=>1162.93260595392,
381=>1163.892761586847,
382=>1164.8519428144,
383=>1165.81014737843,
384=>1166.767373023088,
385=>1167.7236174948296,
386=>1168.6788785424196,
387=>1169.633153916939,
388=>1170.5864413717884,
389=>1171.538738662695,
390=>1172.4900435477166,
391=>1173.4403537872472,
392=>1174.3896671440232,
393=>1175.337981383127,
394=>1176.2852942719942,
395=>1177.2316035804165,
396=>1178.1769070805494,
397=>1179.1212025469158,
398=>1180.0644877564123,
399=>1181.006760488313,
400=>1181.948018524276,
401=>1182.8882596483488,
402=>1183.827481646972,
403=>1184.7656823089867,
404=>1185.7028594256371,
405=>1186.6390107905781,
406=>1187.5741341998787,
407=>1188.5082274520287,
408=>1189.4412883479429,
409=>1190.3733146909663,
410=>1191.3043042868792,
411=>1192.2342549439036,
412=>1193.1631644727067,
413=>1194.091030686407,
414=>1195.0178514005795,
415=>1195.9436244332599,
416=>1196.8683476049505,
417=>1197.792018738626,
418=>1198.7146356597368,
419=>1199.6361961962166,
420=>1200.556698178484,
421=>1201.476139439452,
422=>1202.394517814529,
423=>1203.3118311416267,
424=>1204.228077261164,
425=>1205.1432540160718,
426=>1206.057359251799,
427=>1206.970390816317,
428=>1207.882346560125,
429=>1208.7932243362548,
430=>1209.703022000276,
431=>1210.6117374103012,
432=>1211.519368426991,
433=>1212.425912913558,
434=>1213.3313687357743,
435=>1214.2357337619737,
436=>1215.1390058630584,
437=>1216.0411829125042,
438=>1216.9422627863637,
439=>1217.8422433632738,
440=>1218.7411225244587,
441=>1219.6388981537352,
442=>1220.5355681375195,
443=>1221.4311303648292,
444=>1222.3255827272908,
445=>1223.2189231191435,
446=>1224.111149437244,
447=>1225.0022595810722,
448=>1225.8922514527358,
449=>1226.7811229569747,
450=>1227.6688720011668,
451=>1228.5554964953326,
452=>1229.44099435214,
453=>1230.325363486909,
454=>1231.2086018176174,
455=>1232.0907072649045,
456=>1232.9716777520773,
457=>1233.8515112051145,
458=>1234.730205552672,
459=>1235.6077587260868,
460=>1236.4841686593832,
461=>1237.3594332892762,
462=>1238.2335505551778,
463=>1239.106518399201,
464=>1239.9783347661646,
465=>1240.8489976035985,
466=>1241.7185048617482,
467=>1242.5868544935797,
468=>1243.4540444547845,
469=>1244.3200727037838,
470=>1245.1849372017343,
471=>1246.0486359125323,
472=>1246.9111668028183,
473=>1247.7725278419828,
474=>1248.6327170021696,
475=>1249.491732258282,
476=>1250.349571587987,
477=>1251.2062329717194,
478=>1252.061714392688,
479=>1252.9160138368784,
480=>1253.7691292930604,
481=>1254.6210587527896,
482=>1255.471800210415,
483=>1256.3213516630822,
484=>1257.1697111107374,
485=>1258.0168765561339,
486=>1258.8628460048362,
487=>1259.7076174652238,
488=>1260.5511889484972,
489=>1261.3935584686815,
490=>1262.2347240426311,
491=>1263.0746836900362,
492=>1263.9134354334246,
493=>1264.7509772981684,
494=>1265.5873073124885,
495=>1266.4224235074578,
496=>1267.2563239170074,
497=>1268.0890065779308,
498=>1268.9204695298881,
499=>1269.750710815411,
500=>1270.5797284799073,
501=>1271.4075205716654,
502=>1272.234085141859,
503=>1273.0594202445523,
504=>1273.8835239367027,
505=>1274.7063942781679,
506=>1275.5280293317087,
507=>1276.3484271629936,
508=>1277.1675858406047,
509=>1277.9855034360407,
510=>1278.802178023723,
511=>1279.617607680998,
512=>1280.431790488144,
513=>1281.2447245283745,
514=>1282.0564078878426,
515=>1282.866838655646,
516=>1283.6760149238316,
517=>1284.483934787399,
518=>1285.2905963443063,
519=>1286.095997695474,
520=>1286.9001369447888,
521=>1287.7030121991093,
522=>1288.5046215682696,
523=>1289.3049631650842,
524=>1290.104035105352,
525=>1290.9018355078608,
526=>1291.6983624943928,
527=>1292.493614189727,
528=>1293.2875887216455,
529=>1294.080284220937,
530=>1294.8716988214014,
531=>1295.6618306598539,
532=>1296.4506778761295,
533=>1297.2382386130882,
534=>1298.0245110166181,
535=>1298.8094932356407,
536=>1299.5931834221146,
537=>1300.3755797310407,
538=>1301.156680320465,
539=>1301.936483351485,
540=>1302.7149869882526,
541=>1303.4921893979786,
542=>1304.268088750937,
543=>1305.0426832204703,
544=>1305.8159709829924,
545=>1306.587950217994,
546=>1307.3586191080456,
547=>1308.1279758388034,
548=>1308.8960185990122,
549=>1309.6627455805105,
550=>1310.4281549782345,
551=>1311.192244990222,
552=>1311.955013817617,
553=>1312.7164596646746,
554=>1313.4765807387635,
555=>1314.2353752503718,
556=>1314.9928414131107,
557=>1315.7489774437186,
558=>1316.5037815620647,
559=>1317.257251991155,
560=>1318.0093869571347,
561=>1318.760184689293,
562=>1319.5096434200673,
563=>1320.2577613850476,
564=>1321.0045368229798,
565=>1321.749967975771,
566=>1322.4940530884928,
567=>1323.2367904093862,
568=>1323.9781781898646,
569=>1324.7182146845184,
570=>1325.4568981511202,
571=>1326.1942268506273,
572=>1326.9301990471865,
573=>1327.664813008138,
574=>1328.3980670040203,
575=>1329.1299593085728,
576=>1329.8604881987408,
577=>1330.58965195468,
578=>1331.3174488597592,
579=>1332.043877200566,
580=>1332.7689352669086,
581=>1333.4926213518224,
582=>1334.2149337515725,
583=>1334.9358707656575,
584=>1335.6554306968144,
585=>1336.3736118510224,
586=>1337.090412537506,
587=>1337.8058310687402,
588=>1338.5198657604537,
589=>1339.2325149316337,
590=>1339.943776904528,
591=>1340.6536500046516,
592=>1341.3621325607883,
593=>1342.0692229049957,
594=>1342.7749193726095,
595=>1343.4792203022464,
596=>1344.182124035809,
597=>1344.8836289184887,
598=>1345.5837332987708,
599=>1346.2824355284372,
600=>1346.979733962571,
601=>1347.6756269595598,
602=>1348.3701128811008,
603=>1349.0631900922033,
604=>1349.7548569611927,
605=>1350.4451118597153,
606=>1351.1339531627414,
607=>1351.8213792485685,
608=>1352.5073884988271,
609=>1353.1919792984827,
610=>1353.8751500358399,
611=>1354.5568991025466,
612=>1355.237224893598,
613=>1355.91612580734,
614=>1356.5936002454723,
615=>1357.2696466130542,
616=>1357.9442633185056,
617=>1358.617448773613,
618=>1359.2892013935325,
619=>1359.959519596793,
620=>1360.6284018053002,
621=>1361.2958464443416,
622=>1361.9618519425876,
623=>1362.6264167320978,
624=>1363.2895392483235,
625=>1363.9512179301105,
626=>1364.611451219705,
627=>1365.270237562755,
628=>1365.9275754083155,
629=>1366.5834632088518,
630=>1367.2378994202422,
631=>1367.8908825017834,
632=>1368.5424109161922,
633=>1369.1924831296105,
634=>1369.8410976116088,
635=>1370.4882528351882,
636=>1371.133947276787,
637=>1371.7781794162813,
638=>1372.42094773699,
639=>1373.0622507256785,
640=>1373.7020868725622,
641=>1374.3404546713086,
642=>1374.9773526190434,
643=>1375.6127792163525,
644=>1376.2467329672845,
645=>1376.8792123793569,
646=>1377.5102159635576,
647=>1378.1397422343484,
648=>1378.7677897096705,
649=>1379.394356910945,
650=>1380.0194423630785,
651=>1380.6430445944666,
652=>1381.2651621369957,
653=>1381.8857935260485,
654=>1382.5049373005058,
655=>1383.1225920027512,
656=>1383.7387561786732,
657=>1384.3534283776698,
658=>1384.9666071526515,
659=>1385.5782910600446,
660=>1386.188478659795,
661=>1386.7971685153707,
662=>1387.404359193766,
663=>1388.0100492655047,
664=>1388.6142373046437,
665=>1389.2169218887752,
666=>1389.8181015990317,
667=>1390.4177750200888,
668=>1391.0159407401666,
669=>1391.612597351037,
670=>1392.207743448023,
671=>1392.801377630004,
672=>1393.3934984994198,
673=>1393.9841046622719,
674=>1394.5731947281283,
675=>1395.1607673101255,
676=>1395.7468210249735,
677=>1396.3313544929579,
678=>1396.9143663379427,
679=>1397.495855187375,
680=>1398.0758196722866,
681=>1398.6542584272988,
682=>1399.2311700906243,
683=>1399.806553304071,
684=>1400.3804067130457,
685=>1400.9527289665557,
686=>1401.5235187172143,
687=>1402.0927746212415,
688=>1402.6604953384694,
689=>1403.226679532343,
690=>1403.7913258699261,
691=>1404.354433021902,
692=>1404.915999662578,
693=>1405.4760244698887,
694=>1406.0345061253965,
695=>1406.5914433142998,
696=>1407.1468347254304,
697=>1407.7006790512605,
698=>1408.2529749879047,
699=>1408.8037212351223,
700=>1409.352916496321,
701=>1409.9005594785601,
702=>1410.4466488925536,
703=>1410.9911834526722,
704=>1411.534161876948,
705=>1412.075582887076,
706=>1412.6154452084181,
707=>1413.1537475700056,
708=>1413.690488704542,
709=>1414.2256673484071,
710=>1414.7592822416586,
711=>1415.2913321280357,
712=>1415.8218157549618,
713=>1416.3507318735487,
714=>1416.878079238597,
715=>1417.4038566086015,
716=>1417.9280627457529,
717=>1418.4506964159414,
718=>1418.9717563887582,
719=>1419.4912414375003,
720=>1420.0091503391723,
721=>1420.5254818744888,
722=>1421.0402348278785,
723=>1421.5534079874865,
724=>1422.0650001451768,
725=>1422.5750100965354,
726=>1423.0834366408737,
727=>1423.5902785812305,
728=>1424.0955347243753,
729=>1424.5992038808106,
730=>1425.1012848647754,
731=>1425.6017764942476,
732=>1426.100677590947,
733=>1426.5979869803373,
734=>1427.09370349163,
735=>1427.5878259577867,
736=>1428.0803532155214,
737=>1428.5712841053037,
738=>1429.0606174713614,
739=>1429.5483521616839,
740=>1430.0344870280232,
741=>1430.5190209258985,
742=>1431.001952714598,
743=>1431.4832812571813,
744=>1431.9630054204822,
745=>1432.4411240751128,
746=>1432.9176360954634,
747=>1433.3925403597082,
748=>1433.8658357498052,
749=>1434.3375211515008,
750=>1434.8075954543317,
751=>1435.2760575516272,
752=>1435.7429063405123,
753=>1436.20814072191,
754=>1436.6717596005442,
755=>1437.1337618849423,
756=>1437.5941464874368,
757=>1438.0529123241695,
758=>1438.5100583150925,
759=>1438.9655833839715,
760=>1439.419486458389,
761=>1439.8717664697451,
762=>1440.3224223532616,
763=>1440.7714530479834,
764=>1441.2188574967822,
765=>1441.6646346463576,
766=>1442.1087834472407,
767=>1442.5513028537957,
768=>1442.9921918242235,
769=>1443.4314493205625,
770=>1443.8690743086927,
771=>1444.3050657583372,
772=>1444.7394226430652,
773=>1445.1721439402932,
774=>1445.6032286312893,
775=>1446.0326757011737,
776=>1446.4604841389228,
777=>1446.88665293737,
778=>1447.3111810932091,
779=>1447.7340676069964,
780=>1448.1553114831531,
781=>1448.5749117299677,
782=>1448.9928673595975,
783=>1449.4091773880725,
784=>1449.8238408352963,
785=>1450.2368567250496,
786=>1450.648224084991,
787=>1451.0579419466603,
788=>1451.4660093454813,
789=>1451.8724253207629,
790=>1452.2771889157016,
791=>1452.6802991773848,
792=>1453.0817551567911,
793=>1453.4815559087951,
794=>1453.8797004921676,
795=>1454.2761879695774,
796=>1454.671017407596,
797=>1455.0641878766978,
798=>1455.4556984512628,
799=>1455.8455482095787,
800=>1456.2337362338435,
801=>1456.6202616101666,
802=>1457.0051234285727,
803=>1457.388320783002,
804=>1457.7698527713142,
805=>1458.1497184952884,
806=>1458.5279170606277,
807=>1458.9044475769597,
808=>1459.2793091578392,
809=>1459.652500920749,
810=>1460.0240219871043,
811=>1460.3938714822534,
812=>1460.7620485354794,
813=>1461.1285522800029,
814=>1461.493381852984,
815=>1461.856536395524,
816=>1462.2180150526679,
817=>1462.5778169734058,
818=>1462.9359413106758,
819=>1463.292387221365,
820=>1463.6471538663122,
821=>1464.0002404103093,
822=>1464.3516460221035,
823=>1464.7013698743997,
824=>1465.049411143862,
825=>1465.3957690111156,
826=>1465.740442660749,
827=>1466.0834312813154,
828=>1466.4247340653355,
829=>1466.7643502092983,
830=>1467.1022789136637,
831=>1467.4385193828653,
832=>1467.7730708253093,
833=>1468.1059324533799,
834=>1468.4371034834385,
835=>1468.7665831358274,
836=>1469.0943706348705,
837=>1469.4204652088752,
838=>1469.7448660901346,
839=>1470.0675725149295,
840=>1470.3885837235293,
841=>1470.7078989601946,
842=>1471.0255174731792,
843=>1471.3414385147307,
844=>1471.6556613410933,
845=>1471.968185212509,
846=>1472.2790093932201,
847=>1472.5881331514697,
848=>1472.8955557595045,
849=>1473.2012764935762,
850=>1473.5052946339429,
851=>1473.8076094648713,
852=>1474.1082202746375,
853=>1474.4071263555297,
854=>1474.70432700385,
855=>1474.9998215199146,
856=>1475.2936092080568,
857=>1475.5856893766281,
858=>1475.8760613379998,
859=>1476.1647244085652,
860=>1476.45167790874,
861=>1476.7369211629655,
862=>1477.0204534997085,
863=>1477.3022742514645,
864=>1477.5823827547579,
865=>1477.8607783501445,
866=>1478.1374603822126,
867=>1478.4124281995844,
868=>1478.6856811549183,
869=>1478.9572186049095,
870=>1479.2270399102918,
871=>1479.49514443584,
872=>1479.76153155037,
873=>1480.0262006267403,
874=>1480.2891510418558,
875=>1480.550382176666,
876=>1480.8098934161685,
877=>1481.06768414941,
878=>1481.3237537694881,
879=>1481.5781016735514,
880=>1481.8307272628026,
881=>1482.0816299424991,
882=>1482.3308091219542,
883=>1482.5782642145384,
884=>1482.823994637682,
885=>1483.0679998128749,
886=>1483.310279165669,
887=>1483.5508321256793,
888=>1483.7896581265845,
889=>1484.0267566061298,
890=>1484.262127006127,
891=>1484.4957687724561,
892=>1484.727681355067,
893=>1484.9578642079807,
894=>1485.1863167892898,
895=>1485.4130385611609,
896=>1485.638028989835,
897=>1485.8612875456295,
898=>1486.0828137029387,
899=>1486.3026069402354,
900=>1486.5206667400726,
901=>1486.736992589084,
902=>1486.9515839779847,
903=>1487.1644404015742,
904=>1487.375561358736,
905=>1487.5849463524396,
906=>1487.792594889741,
907=>1487.9985064817847,
908=>1488.202680643804,
909=>1488.4051168951228,
910=>1488.6058147591561,
911=>1488.804773763412,
912=>1489.001993439492,
913=>1489.1974733230927,
914=>1489.3912129540058,
915=>1489.5832118761214,
916=>1489.773469637426,
917=>1489.961985790006,
918=>1490.148759890049,
919=>1490.333791497842,
920=>1490.5170801777751,
921=>1490.6986254983417,
922=>1490.8784270321398,
923=>1491.056484355872,
924=>1491.2327970503477,
925=>1491.4073647004834,
926=>1491.5801868953042,
927=>1491.7512632279436,
928=>1491.920593295646,
929=>1492.0881766997672,
930=>1492.2540130457742,
931=>1492.4181019432476,
932=>1492.580443005882,
933=>1492.7410358514858,
934=>1492.8998801019848,
935=>1493.0569753834202,
936=>1493.212321325951,
937=>1493.365917563855,
938=>1493.5177637355282,
939=>1493.667859483488,
940=>1493.8162044543722,
941=>1493.9627982989396,
942=>1494.1076406720722,
943=>1494.2507312327762,
944=>1494.392069644181,
945=>1494.5316555735403,
946=>1494.6694886922357,
947=>1494.8055686757734,
948=>1494.9398952037882,
949=>1495.0724679600416,
950=>1495.2032866324255,
951=>1495.3323509129602,
952=>1495.4596604977967,
953=>1495.585215087217,
954=>1495.7090143856344,
955=>1495.831058101595,
956=>1495.9513459477785,
957=>1496.0698776409968,
958=>1496.1866529021977,
959=>1496.3016714564633,
960=>1496.4149330330115,
961=>1496.5264373651971,
962=>1496.6361841905114,
963=>1496.7441732505831,
964=>1496.8504042911795,
965=>1496.9548770622064,
966=>1497.0575913177097,
967=>1497.1585468158744,
968=>1497.2577433190263,
969=>1497.3551805936331,
970=>1497.4508584103028,
971=>1497.5447765437862,
972=>1497.6369347729776,
973=>1497.7273328809133,
974=>1497.8159706547742,
975=>1497.902847885885,
976=>1497.9879643697154,
977=>1498.0713199058805,
978=>1498.1529142981403,
979=>1498.2327473544021,
980=>1498.3108188867188,
981=>1498.387128711291,
982=>1498.461676648467,
983=>1498.5344625227417,
984=>1498.60548616276,
985=>1498.6747474013146,
986=>1498.7422460753473,
987=>1498.80798202595,
988=>1498.8719550983637,
989=>1498.9341651419804,
990=>1498.994612010342,
991=>1499.053295561142,
992=>1499.110215656225,
993=>1499.1653721615864,
994=>1499.218764947375,
995=>1499.2703938878908,
996=>1499.3202588615864,
997=>1499.3683597510671,
998=>1499.4146964430925,
999=>1499.4592688285738,
1000=>1499.5020768025772,
1001=>1499.5431202643217,
1002=>1499.5823991171815,
1003=>1499.6199132686838,
1004=>1499.6556626305114,
1005=>1499.6896471185016,
1006=>1499.7218666526464,
1007=>1499.7523211570933,
1008=>1499.7810105601448,
1009=>1499.8079347942587,
1010=>1499.833093796049,
1011=>1499.8564875062857,
1012=>1499.8781158698932,
1013=>1499.8979788359538,
1014=>1499.9160763577052,
1015=>1499.9324083925408,
1016=>1499.9469749020113,
1017=>1499.9597758518237,
1018=>1499.9708112118415,
1019=>1499.980080956084,
1020=>1499.9875850627288,
1021=>1499.993323514109,
1022=>1499.997296296715,
1023=>1499.999503401194,
1024=>1499.9999448223493,
1025=>1499.9986205591426,
1026=>1499.9955306146908,
1027=>1499.9906749962688,
1028=>1499.9840537153077,
1029=>1499.975666787396,
1030=>1499.965514232278,
1031=>1499.9535960738558,
1032=>1499.9399123401874,
1033=>1499.9244630634878,
1034=>1499.9072482801284,
1035=>1499.888268030637,
1036=>1499.867522359698,
1037=>1499.8450113161512,
1038=>1499.820734952994,
1039=>1499.794693327378,
1040=>1499.7668865006121,
1041=>1499.7373145381607,
1042=>1499.705977509643,
1043=>1499.672875488834,
1044=>1499.6380085536643,
1045=>1499.6013767862194,
1046=>1499.562980272739,
1047=>1499.5228191036183,
1048=>1499.4808933734066,
1049=>1499.437203180807,
1050=>1499.3917486286773,
1051=>1499.3445298240285,
1052=>1499.2955468780256,
1053=>1499.244799905986,
1054=>1499.1922890273809,
1055=>1499.138014365834,
1056=>1499.0819760491208,
1057=>1499.0241742091694,
1058=>1498.9646089820596,
1059=>1498.9032805080228,
1060=>1498.840188931441,
1061=>1498.7753344008472,
1062=>1498.7087170689254,
1063=>1498.6403370925086,
1064=>1498.5701946325808,
1065=>1498.498289854274,
1066=>1498.4246229268697,
1067=>1498.3491940237986,
1068=>1498.2720033226383,
1069=>1498.1930510051147,
1070=>1498.1123372571014,
1071=>1498.0298622686182,
1072=>1497.9456262338317,
1073=>1497.8596293510536,
1074=>1497.7718718227425,
1075=>1497.6823538555009,
1076=>1497.5910756600758,
1077=>1497.4980374513589,
1078=>1497.4032394483852,
1079=>1497.3066818743318,
1080=>1497.2083649565197,
1081=>1497.108288926411,
1082=>1497.006454019609,
1083=>1496.9028604758582,
1084=>1496.7975085390435,
1085=>1496.690398457189,
1086=>1496.5815304824582,
1087=>1496.4709048711534,
1088=>1496.3585218837143,
1089=>1496.2443817847181,
1090=>1496.1284848428786,
1091=>1496.010831331046,
1092=>1495.891421526205,
1093=>1495.7702557094763,
1094=>1495.6473341661135,
1095=>1495.5226571855046,
1096=>1495.3962250611698,
1097=>1495.2680380907614,
1098=>1495.1380965760627,
1099=>1495.0064008229886,
1100=>1494.872951141583,
1101=>1494.737747846019,
1102=>1494.6007912545988,
1103=>1494.4620816897518,
1104=>1494.3216194780343,
1105=>1494.179404950129,
1106=>1494.0354384408442,
1107=>1493.8897202891117,
1108=>1493.7422508379886,
1109=>1493.5930304346543,
1110=>1493.4420594304097,
1111=>1493.2893381806782,
1112=>1493.134867045003,
1113=>1492.9786463870469,
1114=>1492.8206765745922,
1115=>1492.6609579795388,
1116=>1492.499490977903,
1117=>1492.3362759498182,
1118=>1492.1713132795328,
1119=>1492.004603355409,
1120=>1491.8361465699236,
1121=>1491.665943319665,
1122=>1491.4939940053337,
1123=>1491.3202990317404,
1124=>1491.144858807806,
1125=>1490.9676737465597,
1126=>1490.788744265139,
1127=>1490.6080707847882,
1128=>1490.4256537308563,
1129=>1490.2414935327984,
1130=>1490.055590624173,
1131=>1489.867945442641,
1132=>1489.6785584299655,
1133=>1489.4874300320103,
1134=>1489.2945606987382,
1135=>1489.0999508842112,
1136=>1488.9036010465888,
1137=>1488.705511648127,
1138=>1488.5056831551767,
1139=>1488.3041160381833,
1140=>1488.1008107716855,
1141=>1487.8957678343138,
1142=>1487.6889877087897,
1143=>1487.4804708819247,
1144=>1487.2702178446189,
1145=>1487.0582290918587,
1146=>1486.8445051227186,
1147=>1486.6290464403573,
1148=>1486.4118535520176,
1149=>1486.192926969025,
1150=>1485.9722672067858,
1151=>1485.749874784788,
1152=>1485.5257502265981,
1153=>1485.2998940598604,
1154=>1485.072306816296,
1155=>1484.8429890317007,
1156=>1484.6119412459457,
1157=>1484.3791640029735,
1158=>1484.1446578507998,
1159=>1483.9084233415092,
1160=>1483.6704610312563,
1161=>1483.4307714802626,
1162=>1483.1893552528163,
1163=>1482.9462129172705,
1164=>1482.7013450460422,
1165=>1482.4547522156108,
1166=>1482.2064350065161,
1167=>1481.9563940033584,
1168=>1481.704629794795,
1169=>1481.4511429735414,
1170=>1481.1959341363677,
1171=>1480.9390038840984,
1172=>1480.68035282161,
1173=>1480.4199815578315,
1174=>1480.1578907057406,
1175=>1479.8940808823636,
1176=>1479.6285527087734,
1177=>1479.361306810089,
1178=>1479.0923438154732,
1179=>1478.8216643581304,
1180=>1478.5492690753072,
1181=>1478.275158608289,
1182=>1477.999333602399,
1183=>1477.7217947069973,
1184=>1477.442542575479,
1185=>1477.1615778652717,
1186=>1476.8789012378356,
1187=>1476.5945133586615,
1188=>1476.3084148972682,
1189=>1476.0206065272016,
1190=>1475.7310889260336,
1191=>1475.4398627753599,
1192=>1475.1469287607983,
1193=>1474.8522875719877,
1194=>1474.5559399025858,
1195=>1474.257886450268,
1196=>1473.9581279167255,
1197=>1473.6566650076636,
1198=>1473.3534984328,
1199=>1473.0486289058636,
1200=>1472.7420571445923,
1201=>1472.433783870731,
1202=>1472.1238098100312,
1203=>1471.8121356922481,
1204=>1471.4987622511392,
1205=>1471.1836902244625,
1206=>1470.8669203539753,
1207=>1470.5484533854315,
1208=>1470.228290068581,
1209=>1469.906431157167,
1210=>1469.582877408924,
1211=>1469.257629585578,
1212=>1468.9306884528414,
1213=>1468.6020547804148,
1214=>1468.2717293419826,
1215=>1467.9397129152119,
1216=>1467.606006281751,
1217=>1467.2706102272277,
1218=>1466.9335255412468,
1219=>1466.5947530173883,
1220=>1466.2542934532062,
1221=>1465.912147650226,
1222=>1465.5683164139432,
1223=>1465.2228005538211,
1224=>1464.8756008832888,
1225=>1464.52671821974,
1226=>1464.1761533845304,
1227=>1463.8239072029755,
1228=>1463.4699805043497,
1229=>1463.1143741218834,
1230=>1462.7570888927617,
1231=>1462.3981256581214,
1232=>1462.0374852630512,
1233=>1461.6751685565864,
1234=>1461.3111763917098,
1235=>1460.945509625349,
1236=>1460.578169118373,
1237=>1460.209155735592,
1238=>1459.838470345754,
1239=>1459.4661138215438,
1240=>1459.0920870395805,
1241=>1458.7163908804148,
1242=>1458.339026228528,
1243=>1457.9599939723291,
1244=>1457.5792950041537,
1245=>1457.1969302202601,
1246=>1456.8129005208298,
1247=>1456.427206809963,
1248=>1456.0398499956773,
1249=>1455.6508309899064,
1250=>1455.260150708496,
1251=>1454.8678100712045,
1252=>1454.4738100016975,
1253=>1454.0781514275484,
1254=>1453.680835280235,
1255=>1453.281862495137,
1256=>1452.8812340115342,
1257=>1452.478950772605,
1258=>1452.075013725423,
1259=>1451.6694238209557,
1260=>1451.2621820140612,
1261=>1450.8532892634867,
1262=>1450.4427465318665,
1263=>1450.0305547857192,
1264=>1449.6167149954456,
1265=>1449.2012281353263,
1266=>1448.7840951835196,
1267=>1448.365317122059,
1268=>1447.9448949368511,
1269=>1447.5228296176736,
1270=>1447.0991221581712,
1271=>1446.6737735558563,
1272=>1446.2467848121037,
1273=>1445.8181569321498,
1274=>1445.3878909250907,
1275=>1444.9559878038776,
1276=>1444.5224485853173,
1277=>1444.0872742900679,
1278=>1443.650465942636,
1279=>1443.2120245713766,
1280=>1442.7719512084882,
1281=>1442.3302468900115,
1282=>1441.886912655828,
1283=>1441.4419495496545,
1284=>1440.9953586190445,
1285=>1440.5471409153822,
1286=>1440.0972974938827,
1287=>1439.645829413588,
1288=>1439.192737737365,
1289=>1438.738023531903,
1290=>1438.281687867711,
1291=>1437.8237318191157,
1292=>1437.364156464258,
1293=>1436.9029628850913,
1294=>1436.440152167379,
1295=>1435.9757254006909,
1296=>1435.5096836784023,
1297=>1435.04202809769,
1298=>1434.5727597595303,
1299=>1434.101879768696,
1300=>1433.6293892337549,
1301=>1433.1552892670657,
1302=>1432.679580984776,
1303=>1432.2022655068206,
1304=>1431.7233439569175,
1305=>1431.2428174625657,
1306=>1430.7606871550424,
1307=>1430.276954169402,
1308=>1429.7916196444698,
1309=>1429.3046847228434,
1310=>1428.816150550887,
1311=>1428.3260182787303,
1312=>1427.8342890602657,
1313=>1427.3409640531438,
1314=>1426.8460444187735,
1315=>1426.349531322318,
1316=>1425.8514259326903,
1317=>1425.3517294225535,
1318=>1424.8504429683157,
1319=>1424.3475677501292,
1320=>1423.8431049518854,
1321=>1423.337055761214,
1322=>1422.8294213694796,
1323=>1422.3202029717777,
1324=>1421.8094017669346,
1325=>1421.2970189575008,
1326=>1420.7830557497527,
1327=>1420.2675133536852,
1328=>1419.7503929830125,
1329=>1419.231695855163,
1330=>1418.7114231912772,
1331=>1418.1895762162048,
1332=>1417.6661561585024,
1333=>1417.1411642504295,
1334=>1416.6146017279457,
1335=>1416.0864698307091,
1336=>1415.5567698020723,
1337=>1415.0255028890788,
1338=>1414.4926703424624,
1339=>1413.9582734166413,
1340=>1413.4223133697178,
1341=>1412.8847914634734,
1342=>1412.345708963367,
1343=>1411.8050671385313,
1344=>1411.2628672617705,
1345=>1410.719110609556,
1346=>1410.1737984620252,
1347=>1409.6269321029765,
1348=>1409.0785128198684,
1349=>1408.5285419038146,
1350=>1407.9770206495814,
1351=>1407.4239503555864,
1352=>1406.8693323238926,
1353=>1406.3131678602072,
1354=>1405.7554582738783,
1355=>1405.1962048778914,
1356=>1404.6354089888669,
1357=>1404.073071927056,
1358=>1403.5091950163383,
1359=>1402.9437795842186,
1360=>1402.376826961825,
1361=>1401.808338483902,
1362=>1401.2383154888125,
1363=>1400.6667593185302,
1364=>1400.0936713186388,
1365=>1399.5190528383291,
1366=>1398.9429052303938,
1367=>1398.365229851226,
1368=>1397.786028060816,
1369=>1397.2053012227477,
1370=>1396.623050704194,
1371=>1396.0392778759162,
1372=>1395.4539841122591,
1373=>1394.8671707911487,
1374=>1394.2788392940874,
1375=>1393.6889910061523,
1376=>1393.0976273159913,
1377=>1392.5047496158202,
1378=>1391.9103593014188,
1379=>1391.3144577721284,
1380=>1390.7170464308474,
1381=>1390.1181266840294,
1382=>1389.5176999416788,
1383=>1388.9157676173475,
1384=>1388.3123311281324,
1385=>1387.7073918946717,
1386=>1387.1009513411407,
1387=>1386.49301089525,
1388=>1385.883571988241,
1389=>1385.2726360548827,
1390=>1384.6602045334685,
1391=>1384.0462788658126,
1392=>1383.4308604972475,
1393=>1382.8139508766194,
1394=>1382.1955514562849,
1395=>1381.575663692109,
1396=>1380.954289043459,
1397=>1380.3314289732048,
1398=>1379.7070849477113,
1399=>1379.0812584368387,
1400=>1378.4539509139358,
1401=>1377.8251638558395,
1402=>1377.1948987428689,
1403=>1376.563157058823,
1404=>1375.929940290977,
1405=>1375.2952499300793,
1406=>1374.659087470347,
1407=>1374.0214544094633,
1408=>1373.3823522485727,
1409=>1372.7417824922795,
1410=>1372.099746648642,
1411=>1371.4562462291706,
1412=>1370.8112827488237,
1413=>1370.164857726004,
1414=>1369.516972682555,
1415=>1368.8676291437575,
1416=>1368.2168286383258,
1417=>1367.5645726984044,
1418=>1366.9108628595645,
1419=>1366.2557006607994,
1420=>1365.5990876445223,
1421=>1364.941025356562,
1422=>1364.2815153461588,
1423=>1363.6205591659614,
1424=>1362.9581583720233,
1425=>1362.2943145237987,
1426=>1361.6290291841399,
1427=>1360.9623039192916,
1428=>1360.29414029889,
1429=>1359.6245398959554,
1430=>1358.9535042868924,
1431=>1358.2810350514842,
1432=>1357.6071337728886,
1433=>1356.9318020376347,
1434=>1356.2550414356201,
1435=>1355.5768535601053,
1436=>1354.8972400077114,
1437=>1354.2162023784158,
1438=>1353.533742275549,
1439=>1352.8498613057895,
1440=>1352.164561079162,
1441=>1351.477843209031,
1442=>1350.7897093120998,
1443=>1350.1001610084047,
1444=>1349.409199921312,
1445=>1348.7168276775142,
1446=>1348.0230459070258,
1447=>1347.3278562431801,
1448=>1346.6312603226238,
1449=>1345.9332597853158,
1450=>1345.2338562745203,
1451=>1344.533051436806,
1452=>1343.8308469220397,
1453=>1343.1272443833832,
1454=>1342.4222454772903,
1455=>1341.7158518635015,
1456=>1341.0080652050415,
1457=>1340.298887168214,
1458=>1339.5883194225985,
1459=>1338.8763636410463,
1460=>1338.1630214996771,
1461=>1337.4482946778726,
1462=>1336.7321848582765,
1463=>1336.0146937267866,
1464=>1335.2958229725546,
1465=>1334.575574287978,
1466=>1333.8539493687,
1467=>1333.1309499136034,
1468=>1332.4065776248062,
1469=>1331.6808342076592,
1470=>1330.9537213707408,
1471=>1330.225240825854,
1472=>1329.4953942880204,
1473=>1328.7641834754788,
1474=>1328.0316101096794,
1475=>1327.2976759152798,
1476=>1326.5623826201418,
1477=>1325.8257319553263,
1478=>1325.0877256550907,
1479=>1324.3483654568834,
1480=>1323.6076531013398,
1481=>1322.8655903322792,
1482=>1322.1221788967,
1483=>1321.3774205447753,
1484=>1320.6313170298495,
1485=>1319.8838701084342,
1486=>1319.135081540203,
1487=>1318.3849530879884,
1488=>1317.633486517777,
1489=>1316.8806835987066,
1490=>1316.1265461030603,
1491=>1315.3710758062628,
1492=>1314.6142744868773,
1493=>1313.8561439266005,
1494=>1313.0966859102582,
1495=>1312.335902225801,
1496=>1311.5737946643007,
1497=>1310.8103650199469,
1498=>1310.04561509004,
1499=>1309.2795466749894,
1500=>1308.5121615783091,
1501=>1307.7434616066125,
1502=>1306.9734485696076,
1503=>1306.2021242800952,
1504=>1305.4294905539618,
1505=>1304.655549210178,
1506=>1303.880302070792,
1507=>1303.1037509609255,
1508=>1302.3258977087714,
1509=>1301.5467441455876,
1510=>1300.7662921056935,
1511=>1299.9845434264646,
1512=>1299.20149994833,
1513=>1298.4171635147668,
1514=>1297.6315359722953,
1515=>1296.8446191704766,
1516=>1296.0564149619058,
1517=>1295.2669252022101,
1518=>1294.4761517500424,
1519=>1293.684096467078,
1520=>1292.8907612180096,
1521=>1292.0961478705435,
1522=>1291.3002582953955,
1523=>1290.503094366285,
1524=>1289.7046579599323,
1525=>1288.9049509560527,
1526=>1288.1039752373536,
1527=>1287.3017326895288,
1528=>1286.4982252012542,
1529=>1285.6934546641844,
1530=>1284.8874229729472,
1531=>1284.0801320251394,
1532=>1283.2715837213227,
1533=>1282.4617799650186,
1534=>1281.6507226627045,
1535=>1280.8384137238081,
1536=>1280.0248550607052,
1537=>1279.2100485887127,
1538=>1278.3939962260856,
1539=>1277.576699894012,
1540=>1276.7581615166082,
1541=>1275.9383830209151,
1542=>1275.1173663368927,
1543=>1274.2951133974166,
1544=>1273.4716261382723,
1545=>1272.6469064981513,
1546=>1271.8209564186468,
1547=>1270.9937778442481,
1548=>1270.1653727223372,
1549=>1269.3357430031833,
1550=>1268.5048906399395,
1551=>1267.672817588636,
1552=>1266.8395258081778,
1553=>1266.0050172603387,
1554=>1265.1692939097566,
1555=>1264.3323577239303,
1556=>1263.4942106732137,
1557=>1262.6548547308105,
1558=>1261.8142918727715,
1559=>1260.9725240779883,
1560=>1260.1295533281898,
1561=>1259.2853816079357,
1562=>1258.4400109046144,
1563=>1257.5934432084362,
1564=>1256.74568051243,
1565=>1255.8967248124377,
1566=>1255.0465781071098,
1567=>1254.1952423979005,
1568=>1253.3427196890639,
1569=>1252.4890119876472,
1570=>1251.63412130349,
1571=>1250.7780496492142,
1572=>1249.9207990402233,
1573=>1249.062371494696,
1574=>1248.2027690335817,
1575=>1247.3419936805963,
1576=>1246.4800474622168,
1577=>1245.6169324076768,
1578=>1244.7526505489611,
1579=>1243.8872039208018,
1580=>1243.0205945606733,
1581=>1242.152824508787,
1582=>1241.2838958080874,
1583=>1240.4138105042462,
1584=>1239.542570645658,
1585=>1238.6701782834366,
1586=>1237.7966354714074,
1587=>1236.9219442661051,
1588=>1236.0461067267681,
1589=>1235.1691249153337,
1590=>1234.2910008964327,
1591=>1233.4117367373847,
1592=>1232.5313345081945,
1593=>1231.6497962815447,
1594=>1230.7671241327935,
1595=>1229.8833201399682,
1596=>1228.998386383761,
1597=>1228.1123249475236,
1598=>1227.2251379172626,
1599=>1226.3368273816343,
1600=>1225.44739543194,
1601=>1224.5568441621222,
1602=>1223.6651756687568,
1603=>1222.7723920510512,
1604=>1221.8784954108373,
1605=>1220.9834878525683,
1606=>1220.0873714833115,
1607=>1219.1901484127454,
1608=>1218.291820753154,
1609=>1217.3923906194218,
1610=>1216.491860129028,
1611=>1215.5902314020434,
1612=>1214.6875065611239,
1613=>1213.783687731505,
1614=>1212.8787770409995,
1615=>1211.9727766199892,
1616=>1211.0656886014222,
1617=>1210.1575151208067,
1618=>1209.2482583162066,
1619=>1208.3379203282364,
1620=>1207.4265033000547,
1621=>1206.5140093773623,
1622=>1205.6004407083938,
1623=>1204.6857994439151,
1624=>1203.7700877372163,
1625=>1202.8533077441084,
1626=>1201.9354616229164,
1627=>1201.0165515344763,
1628=>1200.0965796421285,
1629=>1199.175548111713,
1630=>1198.2534591115646,
1631=>1197.3303148125076,
1632=>1196.406117387851,
1633=>1195.4808690133827,
1634=>1194.5545718673648,
1635=>1193.6272281305291,
1636=>1192.6988399860704,
1637=>1191.7694096196433,
1638=>1190.8389392193549,
1639=>1189.9074309757616,
1640=>1188.9748870818632,
1641=>1188.0413097330973,
1642=>1187.1067011273344,
1643=>1186.1710634648734,
1644=>1185.2343989484357,
1645=>1184.2967097831593,
1646=>1183.3579981765954,
1647=>1182.4182663387023,
1648=>1181.4775164818398,
1649=>1180.5357508207642,
1650=>1179.5929715726238,
1651=>1178.6491809569534,
1652=>1177.704381195667,
1653=>1176.7585745130566,
1654=>1175.8117631357836,
1655=>1174.8639492928746,
1656=>1173.9151352157169,
1657=>1172.9653231380523,
1658=>1172.0145152959717,
1659=>1171.0627139279109,
1660=>1170.1099212746442,
1661=>1169.15613957928,
1662=>1168.2013710872552,
1663=>1167.2456180463296,
1664=>1166.2888827065813,
1665=>1165.3311673203998,
1666=>1164.3724741424835,
1667=>1163.4128054298315,
1668=>1162.4521634417401,
1669=>1161.490550439797,
1670=>1160.5279686878757,
1671=>1159.564420452131,
1672=>1158.599908000991,
1673=>1157.6344336051566,
1674=>1156.6679995375914,
1675=>1155.700608073519,
1676=>1154.7322614904172,
1677=>1153.7629620680118,
1678=>1152.7927120882723,
1679=>1151.8215138354053,
1680=>1150.849369595851,
1681=>1149.8762816582757,
1682=>1148.9022523135677,
1683=>1147.927283854832,
1684=>1146.9513785773843,
1685=>1145.9745387787452,
1686=>1144.996766758636,
1687=>1144.018064818973,
1688=>1143.038435263861,
1689=>1142.0578803995886,
1690=>1141.0764025346236,
1691=>1140.0940039796064,
1692=>1139.1106870473445,
1693=>1138.1264540528082,
1694=>1137.141307313124,
1695=>1136.155249147569,
1696=>1135.1682818775676,
1697=>1134.1804078266832,
1698=>1133.1916293206143,
1699=>1132.2019486871889,
1700=>1131.2113682563581,
1701=>1130.2198903601927,
1702=>1129.227517332875,
1703=>1128.2342515106957,
1704=>1127.2400952320463,
1705=>1126.2450508374154,
1706=>1125.2491206693826,
1707=>1124.2523070726122,
1708=>1123.2546123938487,
1709=>1122.2560389819107,
1710=>1121.2565891876861,
1711=>1120.256265364125,
1712=>1119.2550698662358,
1713=>1118.2530050510793,
1714=>1117.2500732777623,
1715=>1116.2462769074332,
1716=>1115.2416183032756,
1717=>1114.2360998305026,
1718=>1113.229723856352,
1719=>1112.2224927500808,
1720=>1111.2144088829587,
1721=>1110.205474628263,
1722=>1109.195692361273,
1723=>1108.185064459265,
1724=>1107.1735933015052,
1725=>1106.1612812692456,
1726=>1105.148130745718,
1727=>1104.1341441161278,
1728=>1103.119323767649,
1729=>1102.103672089418,
1730=>1101.0871914725294,
1731=>1100.069884310028,
1732=>1099.0517529969054,
1733=>1098.032799930093,
1734=>1097.0130275084568,
1735=>1095.9924381327926,
1736=>1094.9710342058183,
1737=>1093.9488181321701,
1738=>1092.9257923183961,
1739=>1091.9019591729507,
1740=>1090.877321106189,
1741=>1089.851880530361,
1742=>1088.8256398596063,
1743=>1087.7986015099477,
1744=>1086.770767899286,
1745=>1085.7421414473947,
1746=>1084.7127245759132,
1747=>1083.682519708342,
1748=>1082.651529270037,
1749=>1081.619755688203,
1750=>1080.5872013918897,
1751=>1079.5538688119827,
1752=>1078.5197603812016,
1753=>1077.484878534092,
1754=>1076.4492257070206,
1755=>1075.4128043381686,
1756=>1074.375616867527,
1757=>1073.3376657368904,
1758=>1072.2989533898508,
1759=>1071.2594822717924,
1760=>1070.219254829886,
1761=>1069.1782735130835,
1762=>1068.1365407721105,
1763=>1067.0940590594623,
1764=>1066.0508308293968,
1765=>1065.0068585379304,
1766=>1063.9621446428305,
1767=>1062.9166916036106,
1768=>1061.8705018815244,
1769=>1060.8235779395602,
1770=>1059.7759222424336,
1771=>1058.7275372565846,
1772=>1057.6784254501688,
1773=>1056.6285892930537,
1774=>1055.5780312568122,
1775=>1054.5267538147161,
1776=>1053.4747594417308,
1777=>1052.42205061451,
1778=>1051.3686298113894,
1779=>1050.3144995123807,
1780=>1049.2596621991656,
1781=>1048.2041203550912,
1782=>1047.1478764651624,
1783=>1046.0909330160366,
1784=>1045.0332924960194,
1785=>1043.9749573950564,
1786=>1042.9159302047287,
1787=>1041.856213418247,
1788=>1040.7958095304455,
1789=>1039.7347210377757,
1790=>1038.6729504383006,
1791=>1037.6105002316895,
1792=>1036.5473729192115,
1793=>1035.48357100373,
1794=>1034.4190969896963,
1795=>1033.3539533831445,
1796=>1032.2881426916838,
1797=>1031.221667424495,
1798=>1030.1545300923237,
1799=>1029.0867332074736,
1800=>1028.0182792838007,
1801=>1026.9491708367088,
1802=>1025.8794103831424,
1803=>1024.80900044158,
1804=>1023.7379435320305,
1805=>1022.6662421760252,
1806=>1021.5938988966126,
1807=>1020.5209162183528,
1808=>1019.4472966673106,
1809=>1018.3730427710514,
1810=>1017.2981570586319,
1811=>1016.2226420605981,
1812=>1015.1465003089769,
1813=>1014.0697343372706,
1814=>1012.9923466804513,
1815=>1011.9143398749544,
1816=>1010.8357164586735,
1817=>1009.7564789709528,
1818=>1008.6766299525832,
1819=>1007.5961719457948,
1820=>1006.5151074942517,
1821=>1005.4334391430455,
1822=>1004.3511694386897,
1823=>1003.2683009291129,
1824=>1002.1848361636544,
1825=>1001.1007776930563,
1826=>1000.0161280694597,
1827=>998.9308898463961,
1828=>997.8450655787838,
1829=>996.7586578229193,
1830=>995.6716691364742,
1831=>994.5841020784873,
1832=>993.4959592093588,
1833=>992.4072430908449,
1834=>991.3179562860513,
1835=>990.2281013594265,
1836=>989.1376808767575,
1837=>988.0466974051624,
1838=>986.9551535130844,
1839=>985.8630517702865,
1840=>984.7703947478448,
1841=>983.6771850181431,
1842=>982.5834251548653,
1843=>981.4891177329915,
1844=>980.3942653287908,
1845=>979.2988705198147,
1846=>978.2029358848922,
1847=>977.1064640041232,
1848=>976.0094574588721,
1849=>974.911918831762,
1850=>973.8138507066689,
1851=>972.7152556687153,
1852=>971.6161363042642,
1853=>970.5164952009128,
1854=>969.4163349474874,
1855=>968.315658134035,
1856=>967.2144673518197,
1857=>966.1127651933159,
1858=>965.0105542522012,
1859=>963.9078371233516,
1860=>962.8046164028341,
1861=>961.7008946879022,
1862=>960.5966745769875,
1863=>959.4919586696964,
1864=>958.3867495668015,
1865=>957.2810498702372,
1866=>956.1748621830925,
1867=>955.0681891096053,
1868=>953.9610332551566,
1869=>952.8533972262629,
1870=>951.7452836305723,
1871=>950.6366950768568,
1872=>949.5276341750064,
1873=>948.4181035360234,
1874=>947.3081057720162,
1875=>946.197643496192,
1876=>945.0867193228523,
1877=>943.975335867386,
1878=>942.863495746263,
1879=>941.7512015770287,
1880=>940.638455978297,
1881=>939.5252615697451,
1882=>938.4116209721059,
1883=>937.2975368071635,
1884=>936.1830116977462,
1885=>935.0680482677203,
1886=>933.952649141984,
1887=>932.8368169464611,
1888=>931.720554308095,
1889=>930.6038638548428,
1890=>929.4867482156683,
1891=>928.3692100205366,
1892=>927.2512519004074,
1893=>926.1328764872297,
1894=>925.0140864139335,
1895=>923.8948843144261,
1896=>922.7752728235848,
1897=>921.6552545772503,
1898=>920.534832212221,
1899=>919.4140083662469,
1900=>918.2927856780233,
1901=>917.1711667871836,
1902=>916.0491543342948,
1903=>914.9267509608503,
1904=>913.8039593092637,
1905=>912.680782022863,
1906=>911.5572217458835,
1907=>910.4332811234628,
1908=>909.3089628016331,
1909=>908.1842694273166,
1910=>907.0592036483183,
1911=>905.9337681133195,
1912=>904.8079654718724,
1913=>903.6817983743938,
1914=>902.5552694721573,
1915=>901.4283814172895,
1916=>900.301136862762,
1917=>899.1735384623857,
1918=>898.0455888708047,
1919=>896.9172907434898,
1920=>895.7886467367327,
1921=>894.6596595076384,
1922=>893.5303317141207,
1923=>892.4006660148951,
1924=>891.2706650694728,
1925=>890.1403315381535,
1926=>889.0096680820209,
1927=>887.8786773629349,
1928=>886.7473620435253,
1929=>885.6157247871871,
1930=>884.4837682580726,
1931=>883.3514951210859,
1932=>882.2189080418767,
1933=>881.0860096868337,
1934=>879.9528027230779,
1935=>878.8192898184573,
1936=>877.6854736415402,
1937=>876.5513568616088,
1938=>875.4169421486531,
1939=>874.2822321733643,
1940=>873.1472296071291,
1941=>872.0119371220221,
1942=>870.8763573908014,
1943=>869.7404930869011,
1944=>868.6043468844251,
1945=>867.4679214581412,
1946=>866.3312194834741,
1947=>865.1942436365005,
1948=>864.0569965939403,
1949=>862.9194810331534,
1950=>861.781699632131,
1951=>860.6436550694906,
1952=>859.505350024469,
1953=>858.3667871769161,
1954=>857.2279692072891,
1955=>856.0888987966456,
1956=>854.9495786266375,
1957=>853.8100113795049,
1958=>852.6701997380692,
1959=>851.5301463857279,
1960=>850.3898540064463,
1961=>849.2493252847535,
1962=>848.1085629057345,
1963=>846.9675695550249,
1964=>845.8263479188034,
1965=>844.6849006837867,
1966=>843.5432305372226,
1967=>842.4013401668827,
1968=>841.2592322610584,
1969=>840.1169095085525,
1970=>838.9743745986736,
1971=>837.8316302212303,
1972=>836.688679066524,
1973=>835.5455238253423,
1974=>834.4021671889542,
1975=>833.2586118491025,
1976=>832.1148604979978,
1977=>830.970915828312,
1978=>829.8267805331723,
1979=>828.682457306155,
1980=>827.5379488412777,
1981=>826.3932578329955,
1982=>825.2483869761923,
1983=>824.1033389661757,
1984=>822.9581164986706,
1985=>821.8127222698123,
1986=>820.667158976141,
1987=>819.5214293145937,
1988=>818.3755359825001,
1989=>817.2294816775752,
1990=>816.0832690979126,
1991=>814.9369009419788,
1992=>813.7903799086068,
1993=>812.6437086969883,
1994=>811.4968900066698,
1995=>810.3499265375445,
1996=>809.2028209898468,
1997=>808.0555760641452,
1998=>806.9081944613364,
1999=>805.7606788826395,
2000=>804.6130320295874,
2001=>803.4652566040238,
2002=>802.3173553080942,
2003=>801.1693308442406,
2004=>800.0211859151951,
2005=>798.8729232239733,
2006=>797.7245454738683,
2007=>796.5760553684431,
2008=>795.4274556115264,
2009=>794.2787489072045,
2010=>793.1299379598156,
2011=>791.9810254739432,
2012=>790.8320141544099,
2013=>789.6829067062713,
2014=>788.5337058348084,
2015=>787.3844142455231,
2016=>786.2350346441301,
2017=>785.0855697365525,
2018=>783.9360222289134,
2019=>782.7863948275296,
2020=>781.6366902389075,
2021=>780.4869111697341,
2022=>779.3370603268723,
2023=>778.1871404173539,
2024=>777.0371541483732,
2025=>775.8871042272812,
2026=>774.7369933615774,
2027=>773.5868242589064,
2028=>772.4365996270488,
2029=>771.2863221739166,
2030=>770.1359946075457,
2031=>768.9856196360906,
2032=>767.8351999678163,
2033=>766.684738311094,
2034=>765.5342373743935,
2035=>764.3836998662767,
2036=>763.2331284953924,
2037=>762.0825259704684,
2038=>760.9318950003064,
2039=>759.7812382937741,
2040=>758.6305585598008,
2041=>757.4798585073695,
2042=>756.3291408455113,
2043=>755.1784082832988,
2044=>754.0276635298393,
2045=>752.8769092942694,
2046=>751.7261482857471,
2047=>750.5753832134469,
2048=>749.4246167865532,
2049=>748.2738517142532,
2050=>747.1230907057308,
2051=>745.9723364701609,
2052=>744.8215917167014,
2053=>743.6708591544888,
2054=>742.5201414926307,
2055=>741.3694414401995,
2056=>740.2187617062261,
2057=>739.0681049996938,
2058=>737.9174740295318,
2059=>736.7668715046077,
2060=>735.6163001337234,
2061=>734.4657626256068,
2062=>733.3152616889062,
2063=>732.1648000321838,
2064=>731.0143803639096,
2065=>729.8640053924545,
2066=>728.7136778260837,
2067=>727.5634003729514,
2068=>726.4131757410938,
2069=>725.2630066384227,
2070=>724.112895772719,
2071=>722.9628458516269,
2072=>721.8128595826463,
2073=>720.6629396731279,
2074=>719.5130888302662,
2075=>718.3633097610928,
2076=>717.2136051724705,
2077=>716.0639777710868,
2078=>714.9144302634477,
2079=>713.76496535587,
2080=>712.6155857544774,
2081=>711.4662941651922,
2082=>710.3170932937293,
2083=>709.1679858455904,
2084=>708.018974526057,
2085=>706.870062040185,
2086=>705.721251092796,
2087=>704.5725443884741,
2088=>703.4239446315573,
2089=>702.2754545261322,
2090=>701.1270767760269,
2091=>699.9788140848051,
2092=>698.8306691557599,
2093=>697.6826446919064,
2094=>696.5347433959768,
2095=>695.3869679704131,
2096=>694.2393211173611,
2097=>693.0918055386637,
2098=>691.9444239358553,
2099=>690.7971790101537,
2100=>689.6500734624559,
2101=>688.5031099933308,
2102=>687.3562913030123,
2103=>686.2096200913937,
2104=>685.0630990580213,
2105=>683.9167309020878,
2106=>682.7705183224253,
2107=>681.6244640175004,
2108=>680.4785706854069,
2109=>679.3328410238596,
2110=>678.1872777301878,
2111=>677.0418835013295,
2112=>675.8966610338248,
2113=>674.7516130238076,
2114=>673.6067421670044,
2115=>672.462051158722,
2116=>671.3175426938452,
2117=>670.1732194668275,
2118=>669.0290841716878,
2119=>667.8851395020021,
2120=>666.7413881508974,
2121=>665.5978328110456,
2122=>664.4544761746579,
2123=>663.3113209334762,
2124=>662.1683697787696,
2125=>661.0256254013262,
2126=>659.8830904914474,
2127=>658.7407677389415,
2128=>657.5986598331172,
2129=>656.4567694627776,
2130=>655.3150993162131,
2131=>654.1736520811965,
2132=>653.0324304449749,
2133=>651.8914370942653,
2134=>650.7506747152464,
2135=>649.6101459935536,
2136=>648.4698536142723,
2137=>647.3298002619306,
2138=>646.189988620495,
2139=>645.0504213733623,
2140=>643.9111012033543,
2141=>642.7720307927108,
2142=>641.6332128230841,
2143=>640.4946499755313,
2144=>639.3563449305096,
2145=>638.2183003678691,
2146=>637.0805189668467,
2147=>635.9430034060598,
2148=>634.8057563634998,
2149=>633.6687805165261,
2150=>632.532078541859,
2151=>631.395653115575,
2152=>630.259506913099,
2153=>629.1236426091987,
2154=>627.9880628779781,
2155=>626.8527703928711,
2156=>625.7177678266358,
2157=>624.583057851347,
2158=>623.4486431383913,
2159=>622.31452635846,
2160=>621.180710181543,
2161=>620.0471972769224,
2162=>618.9139903131664,
2163=>617.7810919581235,
2164=>616.6485048789143,
2165=>615.5162317419276,
2166=>614.3842752128131,
2167=>613.2526379564748,
2168=>612.1213226370653,
2169=>610.9903319179792,
2170=>609.8596684618466,
2171=>608.7293349305274,
2172=>607.599333985105,
2173=>606.4696682858795,
2174=>605.3403404923617,
2175=>604.2113532632675,
2176=>603.0827092565103,
2177=>601.9544111291955,
2178=>600.8264615376145,
2179=>599.6988631372382,
2180=>598.5716185827107,
2181=>597.4447305278428,
2182=>596.3182016256063,
2183=>595.1920345281278,
2184=>594.0662318866807,
2185=>592.9407963516819,
2186=>591.8157305726835,
2187=>590.691037198367,
2188=>589.5667188765374,
2189=>588.4427782541168,
2190=>587.3192179771372,
2191=>586.1960406907364,
2192=>585.0732490391499,
2193=>583.9508456657054,
2194=>582.8288332128167,
2195=>581.707214321977,
2196=>580.5859916337533,
2197=>579.4651677877791,
2198=>578.34474542275,
2199=>577.2247271764154,
2200=>576.105115685574,
2201=>574.9859135860667,
2202=>573.8671235127705,
2203=>572.7487480995927,
2204=>571.6307899794637,
2205=>570.5132517843319,
2206=>569.3961361451575,
2207=>568.2794456919052,
2208=>567.1631830535391,
2209=>566.0473508580162,
2210=>564.9319517322801,
2211=>563.8169883022542,
2212=>562.702463192837,
2213=>561.5883790278946,
2214=>560.4747384302555,
2215=>559.3615440217033,
2216=>558.2487984229718,
2217=>557.1365042537375,
2218=>556.0246641326146,
2219=>554.9132806771482,
2220=>553.8023565038086,
2221=>552.6918942279842,
2222=>551.5818964639767,
2223=>550.4723658249941,
2224=>549.3633049231437,
2225=>548.2547163694281,
2226=>547.1466027737375,
2227=>546.038966744844,
2228=>544.9318108903949,
2229=>543.8251378169076,
2230=>542.7189501297632,
2231=>541.613250433199,
2232=>540.5080413303042,
2233=>539.403325423013,
2234=>538.2991053120983,
2235=>537.195383597166,
2236=>536.0921628766489,
2237=>534.9894457477992,
2238=>533.8872348066845,
2239=>532.7855326481807,
2240=>531.6843418659653,
2241=>530.5836650525129,
2242=>529.483504799087,
2243=>528.3838636957357,
2244=>527.2847443312846,
2245=>526.186149293331,
2246=>525.0880811682379,
2247=>523.990542541128,
2248=>522.8935359958768,
2249=>521.7970641151077,
2250=>520.7011294801852,
2251=>519.6057346712091,
2252=>518.5108822670082,
2253=>517.4165748451345,
2254=>516.322814981857,
2255=>515.2296052521551,
2256=>514.1369482297134,
2257=>513.0448464869155,
2258=>511.9533025948375,
2259=>510.8623191232423,
2260=>509.7718986405736,
2261=>508.6820437139489,
2262=>507.592756909155,
2263=>506.50404079064106,
2264=>505.4158979215126,
2265=>504.32833086352565,
2266=>503.2413421770806,
2267=>502.15493442121647,
2268=>501.0691101536037,
2269=>499.98387193054015,
2270=>498.89922230694356,
2271=>497.81516383634573,
2272=>496.7316990708872,
2273=>495.64883056131055,
2274=>494.5665608569548,
2275=>493.4848925057485,
2276=>492.40382805420535,
2277=>491.32337004741703,
2278=>490.2435210290474,
2279=>489.1642835413267,
2280=>488.0856601250458,
2281=>487.00765331954887,
2282=>485.93026566272954,
2283=>484.8534996910233,
2284=>483.777357939402,
2285=>482.7018429413683,
2286=>481.62695722894887,
2287=>480.5527033326895,
2288=>479.47908378164743,
2289=>478.4061011033876,
2290=>477.333757823975,
2291=>476.26205646796967,
2292=>475.1909995584201,
2293=>474.12058961685784,
2294=>473.05082916329144,
2295=>471.9817207161995,
2296=>470.9132667925267,
2297=>469.8454699076764,
2298=>468.77833257550503,
2299=>467.71185730831644,
2300=>466.6460466168558,
2301=>465.58090301030387,
2302=>464.5164289962702,
2303=>463.45262708078866,
2304=>462.3894997683107,
2305=>461.32704956169965,
2306=>460.26527896222444,
2307=>459.20419046955465,
2308=>458.143786581753,
2309=>457.0840697952714,
2310=>456.0250426049438,
2311=>454.9667075039808,
2312=>453.9090669839635,
2313=>452.85212353483786,
2314=>451.79587964490906,
2315=>450.7403378008345,
2316=>449.6855004876195,
2317=>448.63137018861073,
2318=>447.5779493854901,
2319=>446.52524055826945,
2320=>445.4732461852841,
2321=>444.4219687431881,
2322=>443.3714107069464,
2323=>442.3215745498314,
2324=>441.2724627434157,
2325=>440.22407775756653,
2326=>439.17642206044,
2327=>438.1294981184757,
2328=>437.0833083963895,
2329=>436.03785535716963,
2330=>434.99314146206973,
2331=>433.94916917060334,
2332=>432.90594094053796,
2333=>431.86345922788956,
2334=>430.82172648691676,
2335=>429.78074517011413,
2336=>428.740517728208,
2337=>427.7010466101497,
2338=>426.66233426311,
2339=>425.62438313247316,
2340=>424.5871956618315,
2341=>423.5507742929798,
2342=>422.5151214659083,
2343=>421.48023961879886,
2344=>420.4461311880178,
2345=>419.41279860811085,
2346=>418.38024431179707,
2347=>417.34847072996325,
2348=>416.31748029165846,
2349=>415.28727542408734,
2350=>414.25785855260574,
2351=>413.2292321007143,
2352=>412.2013984900526,
2353=>411.17436014039396,
2354=>410.1481194696394,
2355=>409.1226788938115,
2356=>408.0980408270498,
2357=>407.0742076816044,
2358=>406.0511818678303,
2359=>405.02896579418206,
2360=>404.00756186720764,
2361=>402.98697249154355,
2362=>401.96720006990756,
2363=>400.9482470030951,
2364=>399.9301156899724,
2365=>398.912808527471,
2366=>397.89632791058216,
2367=>396.88067623235133,
2368=>395.8658558838727,
2369=>394.85186925428184,
2370=>393.8387187307542,
2371=>392.8264066984947,
2372=>391.8149355407351,
2373=>390.80430763872687,
2374=>389.794525371737,
2375=>388.78559111704124,
2376=>387.77750724991904,
2377=>386.7702761436478,
2378=>385.7639001694976,
2379=>384.75838169672454,
2380=>383.75372309256664,
2381=>382.74992672223743,
2382=>381.74699494892053,
2383=>380.744930133764,
2384=>379.7437346358749,
2385=>378.743410812314,
2386=>377.7439610180891,
2387=>376.7453876061512,
2388=>375.7476929273877,
2389=>374.75087933061724,
2390=>373.7549491625843,
2391=>372.75990476795357,
2392=>371.7657484893044,
2393=>370.7724826671248,
2394=>369.78010963980716,
2395=>368.78863174364164,
2396=>367.7980513128111,
2397=>366.8083706793855,
2398=>365.8195921733169,
2399=>364.8317181224325,
2400=>363.84475085243105,
2401=>362.8586926868764,
2402=>361.87354594719193,
2403=>360.8893129526555,
2404=>359.9059960203936,
2405=>358.9235974653766,
2406=>357.94211960041156,
2407=>356.9615647361393,
2408=>355.98193518102704,
2409=>355.00323324136383,
2410=>354.02546122125483,
2411=>353.0486214226158,
2412=>352.07271614516804,
2413=>351.0977476864324,
2414=>350.12371834172455,
2415=>349.15063040414924,
2416=>348.1784861645948,
2417=>347.20728791172786,
2418=>346.2370379319884,
2419=>345.26773850958295,
2420=>344.2993919264811,
2421=>343.3320004624088,
2422=>342.36556639484365,
2423=>341.40009199900913,
2424=>340.4355795478694,
2425=>339.4720313121244,
2426=>338.5094495602031,
2427=>337.54783655826,
2428=>336.58719457016866,
2429=>335.6275258575167,
2430=>334.66883267960014,
2431=>333.7111172934188,
2432=>332.7543819536705,
2433=>331.79862891274485,
2434=>330.84386042072003,
2435=>329.890078725356,
2436=>328.93728607208936,
2437=>327.9854847040284,
2438=>327.0346768619478,
2439=>326.08486478428324,
2440=>325.13605070712555,
2441=>324.18823686421666,
2442=>323.2414254869435,
2443=>322.29561880433306,
2444=>321.3508190430469,
2445=>320.4070284273763,
2446=>319.464249179236,
2447=>318.52248351816047,
2448=>317.5817336612979,
2449=>316.64200182340466,
2450=>315.70329021684086,
2451=>314.7656010515645,
2452=>313.8289365351267,
2453=>312.89329887266564,
2454=>311.95869026690286,
2455=>311.02511291813687,
2456=>310.0925690242384,
2457=>309.16106078064524,
2458=>308.23059038035683,
2459=>307.3011600139298,
2460=>306.37277186947114,
2461=>305.4454281326353,
2462=>304.51913098661754,
2463=>303.5938826121492,
2464=>302.6696851874925,
2465=>301.7465408884359,
2466=>300.8244518882875,
2467=>299.90342035787194,
2468=>298.98344846552413,
2469=>298.06453837708403,
2470=>297.1466922558921,
2471=>296.22991226278396,
2472=>295.3142005560854,
2473=>294.3995592916065,
2474=>293.48599062263816,
2475=>292.5734966999456,
2476=>291.66207967176416,
2477=>290.75174168379357,
2478=>289.8424848791935,
2479=>288.93431139857825,
2480=>288.0272233800112,
2481=>287.121222959001,
2482=>286.21631226849524,
2483=>285.3124934388766,
2484=>284.40976859795677,
2485=>283.5081398709721,
2486=>282.60760938057865,
2487=>281.70817924684627,
2488=>280.8098515872549,
2489=>279.9126285166889,
2490=>279.01651214743214,
2491=>278.12150458916284,
2492=>277.2276079489493,
2493=>276.3348243312436,
2494=>275.44315583787824,
2495=>274.5526045680602,
2496=>273.66317261836593,
2497=>272.77486208273757,
2498=>271.8876750524765,
2499=>271.0016136162389,
2500=>270.11667986003175,
2501=>269.2328758672065,
2502=>268.35020371845536,
2503=>267.4686654918058,
2504=>266.5882632626152,
2505=>265.7089991035673,
2506=>264.83087508466605,
2507=>263.95389327323164,
2508=>263.0780557338948,
2509=>262.2033645285926,
2510=>261.3298217165636,
2511=>260.45742935434174,
2512=>259.58618949575384,
2513=>258.71610419191256,
2514=>257.8471754912129,
2515=>256.9794054393267,
2516=>256.11279607919835,
2517=>255.24734945103904,
2518=>254.38306759232324,
2519=>253.519952537783,
2520=>252.6580063194035,
2521=>251.79723096641823,
2522=>250.93762850530408,
2523=>250.07920095977693,
2524=>249.22195035078585,
2525=>248.36587869650992,
2526=>247.51098801235247,
2527=>246.65728031093641,
2528=>245.8047576020997,
2529=>244.95342189289045,
2530=>244.1032751875626,
2531=>243.25431948757017,
2532=>242.4065567915639,
2533=>241.5599890953858,
2534=>240.71461839206438,
2535=>239.87044667181038,
2536=>239.02747592201172,
2537=>238.18570812722857,
2538=>237.34514526918963,
2539=>236.5057893267866,
2540=>235.66764227606973,
2541=>234.83070609024355,
2542=>233.99498273966162,
2543=>233.16047419182246,
2544=>232.3271824113641,
2545=>231.4951093600606,
2546=>230.66425699681656,
2547=>229.8346272776629,
2548=>229.00622215575197,
2549=>228.1790435813533,
2550=>227.3530935018489,
2551=>226.5283738617279,
2552=>225.70488660258354,
2553=>224.8826336631073,
2554=>224.0616169790851,
2555=>223.24183848339192,
2556=>222.42330010598812,
2557=>221.6060037739145,
2558=>220.78995141128735,
2559=>219.97514493929486,
2560=>219.161586276192,
2561=>218.3492773372958,
2562=>217.53822003498135,
2563=>216.7284162786774,
2564=>215.9198679748606,
2565=>215.1125770270529,
2566=>214.30654533581583,
2567=>213.50177479874606,
2568=>212.69826731047158,
2569=>211.89602476264645,
2570=>211.09504904394748,
2571=>210.2953420400679,
2572=>209.49690563371507,
2573=>208.69974170460455,
2574=>207.90385212945637,
2575=>207.10923878199048,
2576=>206.31590353292222,
2577=>205.52384824995772,
2578=>204.73307479778998,
2579=>203.94358503809428,
2580=>203.15538082952366,
2581=>202.36846402770482,
2582=>201.58283648523332,
2583=>200.7985000516702,
2584=>200.0154565735354,
2585=>199.2337078943067,
2586=>198.45325585441242,
2587=>197.67410229122868,
2588=>196.89624903907463,
2589=>196.11969792920843,
2590=>195.3444507898223,
2591=>194.5705094460384,
2592=>193.79787571990528,
2593=>193.02655143039271,
2594=>192.25653839338793,
2595=>191.48783842169098,
2596=>190.72045332501068,
2597=>189.95438490996048,
2598=>189.1896349800536,
2599=>188.4262053356996,
2600=>187.6640977741995,
2601=>186.90331408974225,
2602=>186.14385607339977,
2603=>185.38572551312302,
2604=>184.6289241937377,
2605=>183.8734538969402,
2606=>183.11931640129364,
2607=>182.36651348222335,
2608=>181.6150469120122,
2609=>180.86491845979754,
2610=>180.11612989156617,
2611=>179.36868297015076,
2612=>178.62257945522504,
2613=>177.87782110330033,
2614=>177.134409667721,
2615=>176.39234689866032,
2616=>175.65163454311676,
2617=>174.9122743449093,
2618=>174.17426804467368,
2619=>173.43761737985847,
2620=>172.70232408472077,
2621=>171.96838989032108,
2622=>171.2358165245215,
2623=>170.50460571197993,
2624=>169.77475917414642,
2625=>169.04627862925895,
2626=>168.31916579234064,
2627=>167.59342237519365,
2628=>166.86905008639644,
2629=>166.14605063129966,
2630=>165.42442571202173,
2631=>164.70417702744578,
2632=>163.9853062732135,
2633=>163.26781514172387,
2634=>162.55170532212753,
2635=>161.83697850032308,
2636=>161.12363635895338,
2637=>160.4116805774014,
2638=>159.70111283178596,
2639=>158.9919347949584,
2640=>158.2841481364984,
2641=>157.5777545227096,
2642=>156.8727556166166,
2643=>156.16915307796012,
2644=>155.46694856319402,
2645=>154.76614372547965,
2646=>154.0667402146844,
2647=>153.3687396773762,
2648=>152.67214375682,
2649=>151.97695409297398,
2650=>151.2831723224856,
2651=>150.59080007868783,
2652=>149.89983899159517,
2653=>149.21029068790017,
2654=>148.5221567909689,
2655=>147.835438920838,
2656=>147.15013869421023,
2657=>146.46625772445088,
2658=>145.78379762158443,
2659=>145.10275999228895,
2660=>144.42314643989505,
2661=>143.74495856438023,
2662=>143.0681979623654,
2663=>142.39286622711154,
2664=>141.71896494851592,
2665=>141.04649571310767,
2666=>140.3754601040448,
2667=>139.7058597011104,
2668=>139.03769608070832,
2669=>138.37097081586012,
2670=>137.7056854762012,
2671=>137.04184162797708,
2672=>136.37944083403897,
2673=>135.71848465384153,
2674=>135.0589746434382,
2675=>134.40091235547777,
2676=>133.74429933920078,
2677=>133.0891371404357,
2678=>132.4354273015956,
2679=>131.78317136167425,
2680=>131.13237085624257,
2681=>130.4830273174449,
2682=>129.83514227399587,
2683=>129.18871725117617,
2684=>128.54375377082977,
2685=>127.9002533513584,
2686=>127.25821750772081,
2687=>126.6176477514274,
2688=>125.9785455905369,
2689=>125.340912529653,
2690=>124.70475006992069,
2691=>124.0700597090231,
2692=>123.43684294117725,
2693=>122.80510125713124,
2694=>122.17483614416051,
2695=>121.54604908606404,
2696=>120.91874156316135,
2697=>120.29291505228844,
2698=>119.66857102679546,
2699=>119.04571095654103,
2700=>118.4243363078914,
2701=>117.80444854371524,
2702=>117.18604912338083,
2703=>116.56913950275259,
2704=>115.9537211341875,
2705=>115.33979546653177,
2706=>114.72736394511742,
2707=>114.11642801175901,
2708=>113.50698910474989,
2709=>112.89904865885921,
2710=>112.29260810532833,
2711=>111.6876688718678,
2712=>111.08423238265277,
2713=>110.48230005832147,
2714=>109.88187331597067,
2715=>109.28295356915271,
2716=>108.68554222787168,
2717=>108.0896406985812,
2718=>107.49525038417994,
2719=>106.90237268400892,
2720=>106.31100899384796,
2721=>105.7211607059129,
2722=>105.13282920885138,
2723=>104.54601588774074,
2724=>103.96072212408376,
2725=>103.37694929580641,
2726=>102.79469877725273,
2727=>102.21397193918403,
2728=>101.63477014877412,
2729=>101.05709476960646,
2730=>100.48094716167122,
2731=>99.90632868136129,
2732=>99.3332406814701,
2733=>98.7616845111877,
2734=>98.19166151609795,
2735=>97.6231730381752,
2736=>97.05622041578124,
2737=>96.49080498366197,
2738=>95.92692807294452,
2739=>95.36459101113348,
2740=>94.8037951221088,
2741=>94.24454172612195,
2742=>93.68683213979318,
2743=>93.1306676761078,
2744=>92.57604964441384,
2745=>92.02297935041872,
2746=>91.47145809618576,
2747=>90.92148718013175,
2748=>90.37306789702347,
2749=>89.82620153797495,
2750=>89.28088939044403,
2751=>88.73713273822966,
2752=>88.19493286146871,
2753=>87.65429103663303,
2754=>87.11520853652667,
2755=>86.57768663028219,
2756=>86.0417265833587,
2757=>85.50732965753753,
2758=>84.97449711092099,
2759=>84.44323019792773,
2760=>83.91353016929065,
2761=>83.38539827205409,
2762=>82.85883574957074,
2763=>82.33384384149758,
2764=>81.81042378379516,
2765=>81.28857680872295,
2766=>80.76830414483709,
2767=>80.2496070169874,
2768=>79.73248664631467,
2769=>79.21694425024737,
2770=>78.702981042499,
2771=>78.19059823306554,
2772=>77.67979702822208,
2773=>77.17057863052025,
2774=>76.6629442387856,
2775=>76.15689504811428,
2776=>75.6524322498708,
2777=>75.14955703168414,
2778=>74.64827057744662,
2779=>74.14857406730971,
2780=>73.65046867768217,
2781=>73.15395558122623,
2782=>72.65903594685619,
2783=>72.16571093973448,
2784=>71.67398172126957,
2785=>71.18384944911304,
2786=>70.69531527715662,
2787=>70.20838035553015,
2788=>69.72304583059815,
2789=>69.23931284495757,
2790=>68.75718253743469,
2791=>68.27665604308277,
2792=>67.79773449317952,
2793=>67.32041901522405,
2794=>66.84471073293457,
2795=>66.37061076624514,
2796=>65.89812023130389,
2797=>65.4272402404697,
2798=>64.95797190230985,
2799=>64.49031632159756,
2800=>64.02427459930902,
2801=>63.55984783262113,
2802=>63.09703711490897,
2803=>62.6358435357422,
2804=>62.17626818088445,
2805=>61.71831213228893,
2806=>61.26197646809703,
2807=>60.80726226263505,
2808=>60.354170586412124,
2809=>59.90270250611741,
2810=>59.452859084617785,
2811=>59.004641380955604,
2812=>58.55805045034538,
2813=>58.11308734417207,
2814=>57.66975310998828,
2815=>57.22804879151181,
2816=>56.78797542862367,
2817=>56.34953405736417,
2818=>55.912725709932374,
2819=>55.477551414682694,
2820=>55.04401219612248,
2821=>54.61210907490954,
2822=>54.181843067850195,
2823=>53.753215187896444,
2824=>53.3262264441438,
2825=>52.90087784182879,
2826=>52.47717038232645,
2827=>52.055105063148744,
2828=>51.63468287794092,
2829=>51.21590481648059,
2830=>50.79877186467388,
2831=>50.38328500455452,
2832=>49.96944521428088,
2833=>49.557253468133695,
2834=>49.146710736513455,
2835=>48.73781798593893,
2836=>48.330576179044215,
2837=>47.92498627457678,
2838=>47.521049227395,
2839=>47.11876598846584,
2840=>46.71813750486319,
2841=>46.319164719765126,
2842=>45.921848572451495,
2843=>45.5261899983027,
2844=>45.13218992879581,
2845=>44.739849291504015,
2846=>44.34916901009376,
2847=>43.96015000432271,
2848=>43.572793190037146,
2849=>43.18709947917023,
2850=>42.803069779739985,
2851=>42.42070499584668,
2852=>42.0400060276711,
2853=>41.660973771472186,
2854=>41.28360911958532,
2855=>40.907912960419594,
2856=>40.533886178456214,
2857=>40.16152965424624,
2858=>39.79084426440829,
2859=>39.421830881627216,
2860=>39.05449037465132,
2861=>38.68882360829036,
2862=>38.32483144341393,
2863=>37.962514736949174,
2864=>37.601874341878556,
2865=>37.24291110723857,
2866=>36.885625878116684,
2867=>36.53001949565032,
2868=>36.17609279702458,
2869=>35.82384661546985,
2870=>35.473281780260095,
2871=>35.12439911671129,
2872=>34.77719944617911,
2873=>34.43168358605692,
2874=>34.08785234977415,
2875=>33.74570654679394,
2876=>33.40524698261186,
2877=>33.06647445875342,
2878=>32.729389772772265,
2879=>32.39399371824902,
2880=>32.06028708478823,
2881=>31.72827065801755,
2882=>31.397945219585154,
2883=>31.069311547158577,
2884=>30.742370414422226,
2885=>30.41712259107601,
2886=>30.09356884283318,
2887=>29.771709931418968,
2888=>29.45154661456843,
2889=>29.133079646024726,
2890=>28.816309775537434,
2891=>28.501237748860717,
2892=>28.187864307751738,
2893=>27.87619018996884,
2894=>27.566216129269037,
2895=>27.25794285540792,
2896=>26.951371094136448,
2897=>26.646501567199948,
2898=>26.343334992336395,
2899=>26.041872083274484,
2900=>25.742113549731926,
2901=>25.444060097414194,
2902=>25.147712428012255,
2903=>24.853071239201768,
2904=>24.56013722464013,
2905=>24.26891107396625,
2906=>23.97939347279828,
2907=>23.691585102731892,
2908=>23.405486641338484,
2909=>23.12109876216425,
2910=>22.838422134728376,
2911=>22.557457424521203,
2912=>22.278205293002657,
2913=>22.00066639760098,
2914=>21.72484139171104,
2915=>21.45073092469272,
2916=>21.17833564186958,
2917=>20.9076561845269,
2918=>20.638693189910896,
2919=>20.37144729122656,
2920=>20.10591911763663,
2921=>19.842109294259558,
2922=>19.580018442168466,
2923=>19.319647178389914,
2924=>19.06099611590173,
2925=>18.80406586363233,
2926=>18.548857026458563,
2927=>18.295370205204904,
2928=>18.04360599664176,
2929=>17.793564993483756,
2930=>17.545247784389176,
2931=>17.29865495395768,
2932=>17.0537870827294,
2933=>16.8106447471838,
2934=>16.56922851973752,
2935=>16.329538968743805,
2936=>16.091576658490794,
2937=>15.855342149200283,
2938=>15.620835997026461,
2939=>15.388058754054441,
2940=>15.157010968299232,
2941=>14.927693183704037,
2942=>14.700105940139451,
2943=>14.474249773401766,
2944=>14.250125215211824,
2945=>14.027732793214227,
2946=>13.807073030975175,
2947=>13.588146447982353,
2948=>13.370953559642544,
2949=>13.155494877281285,
2950=>12.941770908141166,
2951=>12.729782155381372,
2952=>12.519529118075184,
2953=>12.311012291210204,
2954=>12.104232165686199,
2955=>11.899189228314526,
2956=>11.695883961816662,
2957=>11.494316844823288,
2958=>11.294488351872928,
2959=>11.09639895341104,
2960=>10.900049115788647,
2961=>10.70543930126189,
2962=>10.512569967989862,
2963=>10.32144157003438,
2964=>10.13205455735897,
2965=>9.944409375827036,
2966=>9.758506467201528,
2967=>9.574346269143803,
2968=>9.39192921521203,
2969=>9.211255734860856,
2970=>9.032326253440147,
2971=>8.855141192193969,
2972=>8.679700968259567,
2973=>8.506005994666339,
2974=>8.334056680334925,
2975=>8.163853430076415,
2976=>7.995396644590869,
2977=>7.828686720467431,
2978=>7.663724050181827,
2979=>7.500509022096935,
2980=>7.3390420204613065,
2981=>7.179323425407688,
2982=>7.021353612953021,
2983=>6.86513295499708,
2984=>6.710661819321899,
2985=>6.557940569590301,
2986=>6.406969565345776,
2987=>6.257749162011351,
2988=>6.110279710888221,
2989=>5.964561559155982,
2990=>5.820595049871031,
2991=>5.678380521965778,
2992=>5.537918310248301,
2993=>5.3992087454013244,
2994=>5.2622521539810805,
2995=>5.127048858417197,
2996=>4.993599177011447,
2997=>4.861903423937179,
2998=>4.731961909238635,
2999=>4.603774938830156,
3000=>4.477342814495273,
3001=>4.352665833886363,
3002=>4.229744290523854,
3003=>4.108578473794978,
3004=>3.989168668954221,
3005=>3.8715151571213937,
3006=>3.75561821528197,
3007=>3.6414781162856116,
3008=>3.5290951288465067,
3009=>3.4184695175415527,
3010=>3.309601542810924,
3011=>3.2024914609564803,
3012=>3.0971395241417667,
3013=>2.9935459803909907,
3014=>2.891711073589022,
3015=>2.7916350434801416,
3016=>2.6933181256680427,
3017=>2.5967605516149206,
3018=>2.5019625486410177,
3019=>2.4089243399241695,
3020=>2.3176461444992356,
3021=>2.228128177257531,
3022=>2.1403706489462593,
3023=>2.0543737661683963,
3024=>1.9701377313816693,
3025=>1.887662742898442,
3026=>1.806948994885147,
3027=>1.7279966773617161,
3028=>1.6508059762014682,
3029=>1.5753770731301984,
3030=>1.501710145726065,
3031=>1.4298053674193625,
3032=>1.3596629074912698,
3033=>1.2912829310746474,
3034=>1.224665599152786,
3035=>1.1598110685590655,
3036=>1.0967194919772965,
3037=>1.0353910179403556,
3038=>0.9758257908306405,
3039=>0.9180239508792738,
3040=>0.8619856341661034,
3041=>0.8077109726191338,
3042=>0.7552000940140715,
3043=>0.7044531219745522,
3044=>0.6554701759715726,
3045=>0.6082513713228082,
3046=>0.5627968191930677,
3047=>0.5191066265934978,
3048=>0.4771808963816966,
3049=>0.43701972726091753,
3050=>0.39862321378063825,
3051=>0.36199144633553715,
3052=>0.3271245111659482,
3053=>0.2940224903570652,
3054=>0.26268546183939634,
3055=>0.23311349938785497,
3056=>0.20530667262210045,
3057=>0.17926504700619716,
3058=>0.15498868384872821,
3059=>0.1324776403021133,
3060=>0.11173196936294971,
3061=>0.09275171987155773,
3062=>0.07553693651220783,
3063=>0.060087659812552374,
3064=>0.046403926144193974,
3065=>0.0344857677220034,
3066=>0.024333212604005894,
3067=>0.01594628469217696,
3068=>0.00932500373107814,
3069=>0.004469385309107565,
3070=>0.0013794408574767658,
3071=>5.517765055174095e-05,
3072=>0.0004965988060803284,
3073=>0.0027037032849648313,
3074=>0.006676485890920958,
3075=>0.012414937271159943,
3076=>0.0199190439159338,
3077=>0.029188788158649004,
3078=>0.04022414817632125,
3079=>0.05302509798855226,
3080=>0.06759160745923509,
3081=>0.08392364229496252,
3082=>0.1020211640461639,
3083=>0.12188413010665045,
3084=>0.143512493714411,
3085=>0.16690620395081623,
3086=>0.19206520574130082,
3087=>0.21898943985524966,
3088=>0.24767884290668007,
3089=>0.27813334735355966,
3090=>0.3103528814983747,
3091=>0.34433736948858495,
3092=>0.38008673131628257,
3093=>0.4176008828186468,
3094=>0.45687973567817153,
3095=>0.4979231974227787,
3096=>0.5407311714260459,
3097=>0.5853035569074336,
3098=>0.6316402489327402,
3099=>0.6797411384137604,
3100=>0.7296061121093089,
3101=>0.7812350526249929,
3102=>0.834627838413553,
3103=>0.8897843437750907,
3104=>0.9467044388578643,
3105=>1.0053879896578337,
3106=>1.0658348580195707,
3107=>1.1280449016361445,
3108=>1.192017974049918,
3109=>1.2577539246525475,
3110=>1.3252525986853243,
3111=>1.3945138372399697,
3112=>1.4655374772581808,
3113=>1.5383233515331085,
3114=>1.6128712887089023,
3115=>1.6891811132811654,
3116=>1.767252645597864,
3117=>1.8470857018595552,
3118=>1.9286800941196134,
3119=>2.0120356302844584,
3120=>2.097152114114806,
3121=>2.1840293452256674,
3122=>2.2726671190865773,
3123=>2.363065227022389,
3124=>2.4552234562136164,
3125=>2.549141589697342,
3126=>2.6448194063669916,
3127=>2.7422566809735827,
3128=>2.841453184125612,
3129=>2.9424086822903064,
3130=>3.045122937793508,
3131=>3.149595708820584,
3132=>3.255826749416883,
3133=>3.3638158094885284,
3134=>3.473562634802761,
3135=>3.585066966988279,
3136=>3.698328543536718,
3137=>3.8133470978024206,
3138=>3.930122359003235,
3139=>4.048654052221764,
3140=>4.16894189840491,
3141=>4.290985614365695,
3142=>4.4147849127832615,
3143=>4.540339502203324,
3144=>4.667649087039763,
3145=>4.796713367574398,
3146=>4.927532039958237,
3147=>5.060104796211931,
3148=>5.194431324226457,
3149=>5.3305113077642545,
3150=>5.468344426459566,
3151=>5.607930355819235,
3152=>5.749268767223725,
3153=>5.892359327927693,
3154=>6.037201701060553,
3155=>6.183795545627959,
3156=>6.332140516511799,
3157=>6.482236264471567,
3158=>6.63408243614515,
3159=>6.787678674048948,
3160=>6.943024616579805,
3161=>7.100119898015237,
3162=>7.258964148514224,
3163=>7.419556994118125,
3164=>7.581898056752266,
3165=>7.745986954225714,
3166=>7.911823300232754,
3167=>8.0794067043538,
3168=>8.248736772056418,
3169=>8.41981310469589,
3170=>8.592635299516473,
3171=>8.767202949652187,
3172=>8.943515644127956,
3173=>9.121572967860175,
3174=>9.301374501658188,
3175=>9.482919822224858,
3176=>9.666208502158042,
3177=>9.851240109950936,
3178=>10.038014209993776,
3179=>10.226530362574067,
3180=>10.416788123878746,
3181=>10.608787045994063,
3182=>10.802526676907405,
3183=>10.99800656050786,
3184=>11.195226236587928,
3185=>11.394185240843854,
3186=>11.594883104877226,
3187=>11.797319356195999,
3188=>12.001493518215284,
3189=>12.207405110258946,
3190=>12.415053647560512,
3191=>12.624438641264078,
3192=>12.835559598425789,
3193=>13.048416022015317,
3194=>13.263007410916202,
3195=>13.47933325992733,
3196=>13.697393059764408,
3197=>13.917186297061335,
3198=>14.13871245437042,
3199=>14.361971010164893,
3200=>14.586961438839012,
3201=>14.81368321071011,
3202=>15.042135792019167,
3203=>15.272318644932852,
3204=>15.504231227543755,
3205=>15.737872993872998,
3206=>15.973243393870234,
3207=>16.210341873415473,
3208=>16.44916787432078,
3209=>16.689720834330956,
3210=>16.932000187124913,
3211=>17.176005362317937,
3212=>17.421735785461465,
3213=>17.66919087804581,
3214=>17.918370057500738,
3215=>18.169272737197275,
3216=>18.421898326448513,
3217=>18.67624623051188,
3218=>18.932315850589816,
3219=>19.190106583831493,
3220=>19.44961782333405,
3221=>19.710848958144197,
3222=>19.973799373259567,
3223=>20.238468449629977,
3224=>20.50485556415981,
3225=>20.772960089707908,
3226=>21.042781395090515,
3227=>21.314318845081743,
3228=>21.587571800415617,
3229=>21.862539617787434,
3230=>22.139221649855358,
3231=>22.417617245242013,
3232=>22.69772574853539,
3233=>22.97954650029135,
3234=>23.263078837034527,
3235=>23.548322091259934,
3236=>23.83527559143488,
3237=>24.123938662,
3238=>24.41431062337176,
3239=>24.706390791943136,
3240=>25.000178480085196,
3241=>25.295672996149847,
3242=>25.592873644470046,
3243=>25.89177972536254,
3244=>26.192390535128766,
3245=>26.49470536605702,
3246=>26.7987235064237,
3247=>27.104444240495354,
3248=>27.41186684853028,
3249=>27.72099060677988,
3250=>28.031814787490703,
3251=>28.344338658906622,
3252=>28.65856148526916,
3253=>28.97448252682068,
3254=>29.292101039805175,
3255=>29.611416276470663,
3256=>29.932427485070434,
3257=>30.255133909865208,
3258=>30.57953479112473,
3259=>30.905629365129357,
3260=>31.233416864172455,
3261=>31.56289651656141,
3262=>31.894067546620136,
3263=>32.226929174690554,
3264=>32.56148061713486,
3265=>32.89772108633622,
3266=>33.235649790701814,
3267=>33.575265934664685,
3268=>33.91656871868463,
3269=>34.25955733925116,
3270=>34.60423098888441,
3271=>34.9505888561381,
3272=>35.298630125600425,
3273=>35.648353977896704,
3274=>35.999759589690825,
3275=>36.35284613368776,
3276=>36.70761277863471,
3277=>37.06405868932404,
3278=>37.4221830265941,
3279=>37.78198494733215,
3280=>38.143463604476096,
3281=>38.50661814701607,
3282=>38.87144771999715,
3283=>39.23795146452062,
3284=>39.60612851774658,
3285=>39.97597801289555,
3286=>40.34749907925118,
3287=>40.72069084216082,
3288=>41.095552423039976,
3289=>41.47208293937206,
3290=>41.85028150471146,
3291=>42.23014722868584,
3292=>42.61167921699791,
3293=>42.99487657142731,
3294=>43.37973838983339,
3295=>43.76626376615661,
3296=>44.15445179042115,
3297=>44.54430154873717,
3298=>44.935812123302185,
3299=>45.32898259240403,
3300=>45.72381203042278,
3301=>46.12029950783244,
3302=>46.51844409120463,
3303=>46.91824484320864,
3304=>47.319700822615346,
3305=>47.72281108429843,
3306=>48.12757467923723,
3307=>48.533990654518675,
3308=>48.94205805333968,
3309=>49.35177591500906,
3310=>49.76314327495038,
3311=>50.17615916470345,
3312=>50.59082261192748,
3313=>51.007132640402574,
3314=>51.425088270032234,
3315=>51.844688516846645,
3316=>52.26593239300348,
3317=>52.68881890679086,
3318=>53.113347062630055,
3319=>53.53951586107712,
3320=>53.967324298826156,
3321=>54.39677136871069,
3322=>54.82785605970673,
3323=>55.26057735693496,
3324=>55.694934241662736,
3325=>56.130925691307425,
3326=>56.568550679437635,
3327=>57.00780817577663,
3328=>57.44869714620404,
3329=>57.89121655275903,
3330=>58.335365353642146,
3331=>58.78114250321755,
3332=>59.22854695201636,
3333=>59.677577646738314,
3334=>60.12823353025476,
3335=>60.58051354161091,
3336=>61.03441661602835,
3337=>61.48994168490765,
3338=>61.94708767583063,
3339=>62.405853512563226,
3340=>62.866238115057854,
3341=>63.32824039945547,
3342=>63.79185927808976,
3343=>64.25709365948751,
3344=>64.72394244837255,
3345=>65.19240454566807,
3346=>65.66247884849895,
3347=>66.13416425019454,
3348=>66.60745964029172,
3349=>67.08236390453635,
3350=>67.55887592488716,
3351=>68.03699457951757,
3352=>68.51671874281874,
3353=>68.99804728540198,
3354=>69.48097907410147,
3355=>69.96551297197652,
3356=>70.45164783831592,
3357=>70.93938252863836,
3358=>71.42871589469621,
3359=>71.91964678447857,
3360=>72.41217404221322,
3361=>72.90629650836979,
3362=>73.40201301966249,
3363=>73.89932240905296,
3364=>74.39822350575218,
3365=>74.8987151352245,
3366=>75.40079611918941,
3367=>75.90446527562472,
3368=>76.40972141876921,
3369=>76.91656335912603,
3370=>77.4249899034644,
3371=>77.9349998548231,
3372=>78.4465920125134,
3373=>78.95976517212125,
3374=>79.47451812551105,
3375=>79.99084966082751,
3376=>80.50875856249934,
3377=>81.02824361124158,
3378=>81.54930358405852,
3379=>82.0719372542469,
3380=>82.59614339139853,
3381=>83.12192076140286,
3382=>83.64926812645115,
3383=>84.17818424503776,
3384=>84.70866787196405,
3385=>85.24071775834113,
3386=>85.77433265159254,
3387=>86.30951129545758,
3388=>86.84625242999425,
3389=>87.38455479158176,
3390=>87.92441711292383,
3391=>88.46583812305187,
3392=>89.00881654732768,
3393=>89.55335110744636,
3394=>90.09944052143987,
3395=>90.64708350367903,
3396=>91.19627876487777,
3397=>91.74702501209526,
3398=>92.29932094873936,
3399=>92.85316527456973,
3400=>93.40855668570032,
3401=>93.96549387460334,
3402=>94.52397553011167,
3403=>95.08400033742191,
3404=>95.64556697809803,
3405=>96.20867413007375,
3406=>96.77332046765684,
3407=>97.33950466153067,
3408=>97.90722537875831,
3409=>98.47648128278558,
3410=>99.04727103344408,
3411=>99.61959328695434,
3412=>100.19344669592897,
3413=>100.76882990937577,
3414=>101.34574157270129,
3415=>101.92418032771343,
3416=>102.5041448126251,
3417=>103.08563366205738,
3418=>103.66864550704224,
3419=>104.25317897502623,
3420=>104.8392326898744,
3421=>105.42680527187167,
3422=>106.0158953377279,
3423=>106.60650150057995,
3424=>107.19862236999575,
3425=>107.79225655197706,
3426=>108.38740264896296,
3427=>108.98405925983332,
3428=>109.58222497991142,
3429=>110.18189840096818,
3430=>110.783078111225,
3431=>111.38576269535668,
3432=>111.98995073449521,
3433=>112.59564080623397,
3434=>113.20283148462931,
3435=>113.81152134020488,
3436=>114.42170893995512,
3437=>115.03339284734841,
3438=>115.64657162233016,
3439=>116.26124382132673,
3440=>116.87740799724872,
3441=>117.49506269949393,
3442=>118.11420647395141,
3443=>118.73483786300426,
3444=>119.35695540553354,
3445=>119.9805576369215,
3446=>120.60564308905487,
3447=>121.23221029032936,
3448=>121.86025776565134,
3449=>122.48978403644242,
3450=>123.120787620643,
3451=>123.75326703271548,
3452=>124.38722078364754,
3453=>125.02264738095641,
3454=>125.65954532869125,
3455=>126.29791312743794,
3456=>126.93774927432139,
3457=>127.57905226301,
3458=>128.2218205837188,
3459=>128.86605272321265,
3460=>129.51174716481148,
3461=>130.15890238839108,
3462=>130.80751687038924,
3463=>131.45758908380765,
3464=>132.1091174982165,
3465=>132.76210057975754,
3466=>133.41653679114813,
3467=>134.07242459168435,
3468=>134.72976243724497,
3469=>135.38854878029497,
3470=>136.0487820698894,
3471=>136.71046075167658,
3472=>137.3735832679016,
3473=>138.03814805741195,
3474=>138.70415355565808,
3475=>139.37159819469946,
3476=>140.04048040320686,
3477=>140.71079860646728,
3478=>141.38255122638668,
3479=>142.0557366814943,
3480=>142.7303533869458,
3481=>143.40639975452757,
3482=>144.08387419266,
3483=>144.76277510640193,
3484=>145.44310089745352,
3485=>146.12484996416026,
3486=>146.80802070151697,
3487=>147.49261150117252,
3488=>148.17862075143114,
3489=>148.86604683725852,
3490=>149.55488814028445,
3491=>150.245143038807,
3492=>150.9368099077965,
3493=>151.62988711889898,
3494=>152.32437304043992,
3495=>153.020266037429,
3496=>153.7175644715628,
3497=>154.41626670122912,
3498=>155.11637108151115,
3499=>155.81787596419065,
3500=>156.52077969775314,
3501=>157.22508062739018,
3502=>157.93077709500392,
3503=>158.6378674392115,
3504=>159.34634999534808,
3505=>160.05622309547152,
3506=>160.767485068366,
3507=>161.48013423954592,
3508=>162.19416893125958,
3509=>162.90958746249385,
3510=>163.62638814897753,
3511=>164.3445693031855,
3512=>165.06412923434243,
3513=>165.78506624842714,
3514=>166.5073786481771,
3515=>167.231064733091,
3516=>167.95612279943373,
3517=>168.68255114024032,
3518=>169.41034804531967,
3519=>170.13951180125878,
3520=>170.87004069142745,
3521=>171.60193299597984,
3522=>172.3351869918621,
3523=>173.06980095281335,
3524=>173.8057731493725,
3525=>174.54310184887947,
3526=>175.28178531548144,
3527=>176.02182181013552,
3528=>176.76320959061377,
3529=>177.50594691150707,
3530=>178.25003202422909,
3531=>178.99546317702038,
3532=>179.7422386149526,
3533=>180.49035657993284,
3534=>181.23981531070706,
3535=>181.99061304286533,
3536=>182.74274800884507,
3537=>183.496218437935,
3538=>184.25102255628133,
3539=>185.0071585868891,
3540=>185.76462474962807,
3541=>186.52341926123643,
3542=>187.28354033532526,
3543=>188.0449861823828,
3544=>188.80775500977802,
3545=>189.5718450217655,
3546=>190.33725441948945,
3547=>191.10398140098778,
3548=>191.8720241611967,
3549=>192.64138089195444,
3550=>193.41204978200585,
3551=>194.18402901700722,
3552=>194.9573167795295,
3553=>195.73191124906293,
3554=>196.50781060202144,
3555=>197.2850130117473,
3556=>198.0635166485149,
3557=>198.84331967953494,
3558=>199.6244202689594,
3559=>200.40681657788537,
3560=>201.19050676435927,
3561=>201.97548898338198,
3562=>202.76176138691199,
3563=>203.5493221238703,
3564=>204.338169340146,
3565=>205.12830117859835,
3566=>205.9197157790627,
3567=>206.71241127835424,
3568=>207.50638581027283,
3569=>208.30163750560712,
3570=>209.09816449213895,
3571=>209.89596489464805,
3572=>210.69503683491575,
3573=>211.4953784317304,
3574=>212.29698780089075,
3575=>213.09986305521124,
3576=>213.9040023045261,
3577=>214.70940365569334,
3578=>215.51606521260067,
3579=>216.32398507616824,
3580=>217.13316134435377,
3581=>217.94359211215726,
3582=>218.7552754716254,
3583=>219.5682095118558,
3584=>220.38239231900184,
3585=>221.19782197627694,
3586=>222.01449656395914,
3587=>222.8324141593954,
3588=>223.65157283700648,
3589=>224.47197066829153,
3590=>225.29360572183168,
3591=>226.1164760632969,
3592=>226.94057975544752,
3593=>227.7659148581406,
3594=>228.5924794283343,
3595=>229.42027152009246,
3596=>230.24928918458875,
3597=>231.07953047011165,
3598=>231.91099342206905,
3599=>232.74367608299247,
3600=>233.5775764925421,
3601=>234.41269268751148,
3602=>235.24902270183145,
3603=>236.08656456657548,
3604=>236.92531630996336,
3605=>237.76527595736832,
3606=>238.6064415313183,
3607=>239.44881105150245,
3608=>240.2923825347758,
3609=>241.13715399516354,
3610=>241.9831234438659,
3611=>242.83028888926253,
3612=>243.67864833691777,
3613=>244.52819978958468,
3614=>245.3789412472102,
3615=>246.2308707069397,
3616=>247.0839861631216,
3617=>247.9382856073118,
3618=>248.79376702828023,
3619=>249.65042841201267,
3620=>250.50826774171753,
3621=>251.3672829978301,
3622=>252.2274721580169,
3623=>253.08883319718132,
3624=>253.95136408746743,
3625=>254.81506279826544,
3626=>255.67992729621602,
3627=>256.5459555452154,
3628=>257.4131455064202,
3629=>258.28149513825167,
3630=>259.1510023964015,
3631=>260.0216652338349,
3632=>260.89348160079857,
3633=>261.7664494448218,
3634=>262.6405667107234,
3635=>263.51583134061656,
3636=>264.3922412739128,
3637=>265.2697944473277,
3638=>266.1484887948851,
3639=>267.0283222479224,
3640=>267.90929273509533,
3641=>268.7913981823825,
3642=>269.6746365130908,
3643=>270.55900564785986,
3644=>271.4445035046667,
3645=>272.3311279988325,
3646=>273.2188770430248,
3647=>274.1077485472638,
3648=>274.9977404189274,
3649=>275.88885056275615,
3650=>276.78107688085674,
3651=>277.6744172727094,
3652=>278.5688696351711,
3653=>279.4644318624809,
3654=>280.36110184626506,
3655=>281.25887747554134,
3656=>282.15775663672605,
3657=>283.0577372136361,
3658=>283.95881708749585,
3659=>284.86099413694143,
3660=>285.7642662380263,
3661=>286.6686312642257,
3662=>287.574087086442,
3663=>288.4806315730092,
3664=>289.3882625896988,
3665=>290.29697799972416,
3666=>291.2067756637455,
3667=>292.1176534398753,
3668=>293.02960918368285,
3669=>293.942640748201,
3670=>294.8567459839282,
3671=>295.77192273883594,
3672=>296.68816885837305,
3673=>297.60548218547086,
3674=>298.523860560548,
3675=>299.4433018215158,
3676=>300.3638038037836,
3677=>301.2853643402631,
3678=>302.2079812613742,
3679=>303.1316523950497,
3680=>304.0563755667404,
3681=>304.98214859942016,
3682=>305.9089693135925,
3683=>306.8368355272929,
3684=>307.76574505609614,
3685=>308.69569571312064,
3686=>309.6266853090338,
3687=>310.558711652057,
3688=>311.49177254797115,
3689=>312.42586580012124,
3690=>313.360989209422,
3691=>314.2971405743629,
3692=>315.2343176910134,
3693=>316.1725183530279,
3694=>317.1117403516514,
3695=>318.0519814757237,
3696=>318.99323951168685,
3697=>319.93551224358754,
3698=>320.87879745308385,
3699=>321.82309291945046,
3700=>322.76839641958344,
3701=>323.7147057280058,
3702=>324.66201861687284,
3703=>325.61033285597676,
3704=>326.55964621275274,
3705=>327.5099564522835,
3706=>328.4612613373051,
3707=>329.4135586282116,
3708=>330.3668460830606,
3709=>331.32112145758,
3710=>332.27638250517015,
3711=>333.23262697691166,
3712=>334.1898526215698,
3713=>335.1480571855999,
3714=>336.10723841315274,
3715=>337.06739404607976,
3716=>338.0285218239384,
3717=>338.9906194839975,
3718=>339.9536847612424,
3719=>340.9177153883806,
3720=>341.88270909584685,
3721=>342.8486636118085,
3722=>343.81557666217066,
3723=>344.7834459705831,
3724=>345.7522692584428,
3725=>346.7220442449015,
3726=>347.6927686468704,
3727=>348.66444017902535,
3728=>349.6370565538125,
3729=>350.6106154814538,
3730=>351.585114669952,
3731=>352.56055182509624,
3732=>353.53692465046754,
3733=>354.514230847444,
3734=>355.49246811520663,
3735=>356.47163415074345,
3736=>357.45172664885814,
3737=>358.4327433021711,
3738=>359.4146818011279,
3739=>360.3975398340038,
3740=>361.38131508690907,
3741=>362.366005243795,
3742=>363.3516079864584,
3743=>364.3381209945483,
3744=>365.32554194557025,
3745=>366.3138685148925,
3746=>367.30309837575106,
3747=>368.29322919925556,
3748=>369.28425865439397,
3749=>370.27618440804025,
3750=>371.2690041249567,
3751=>372.26271546780134,
3752=>373.2573160971333,
3753=>374.252803671418,
3754=>375.24917584703286,
3755=>376.24643027827267,
3756=>377.24456461735514,
3757=>378.2435765144266,
3758=>379.24346361756716,
3759=>380.2442235727967,
3760=>381.2458540240802,
3761=>382.248352613333,
3762=>383.25171698042635,
3763=>384.2559447631948,
3764=>385.26103359743865,
3765=>386.26698111693145,
3766=>387.2737849534253,
3767=>388.2814427366564,
3768=>389.28995209435027,
3769=>390.299310652228,
3770=>391.30951603401104,
3771=>392.32056586142767,
3772=>393.33245775421767,
3773=>394.3451893301387,
3774=>395.35875820497154,
3775=>396.37316199252507,
3776=>397.3883983046451,
3777=>398.40446475121377,
3778=>399.42135894016127,
3779=>400.4390784774686,
3780=>401.4576209671737,
3781=>402.4769840113769,
3782=>403.49716521024686,
3783=>404.51816216202604,
3784=>405.53997246303646,
3785=>406.5625937076855,
3786=>407.58602348847035,
3787=>408.6102593959868,
3788=>409.63529901893116,
3789=>410.6611399441078,
3790=>411.6877797564349,
3791=>412.71521603894985,
3792=>413.7434463728149,
3793=>414.7724683373228,
3794=>415.8022795099028,
3795=>416.8328774661261,
3796=>417.8642597797115,
3797=>418.89642402253145,
3798=>419.9293677646173,
3799=>420.9630885741649,
3800=>421.9975840175423,
3801=>423.03285165929213,
3802=>424.06888906213976,
3803=>425.1056937869983,
3804=>426.14326339297435,
3805=>427.1815954373738,
3806=>428.2206874757077,
3807=>429.2605370616976,
3808=>430.301141747282,
3809=>431.3424990826213,
3810=>432.3846066161043,
3811=>433.4274618943535,
3812=>434.4710624622309,
3813=>435.5154058628437,
3814=>436.56048963755165,
3815=>437.6063113259699,
3816=>438.652868465977,
3817=>439.7001585937199,
3818=>440.74817924362014,
3819=>441.79692794837916,
3820=>442.84640223898464,
3821=>443.8965996447159,
3822=>444.9475176931499,
3823=>445.9991539101671,
3824=>447.051505819957,
3825=>448.10457094502453,
3826=>449.1583468061946,
3827=>450.21283092262087,
3828=>451.2680208117878,
3829=>452.3239139895187,
3830=>453.3805079699814,
3831=>454.4378002656937,
3832=>455.4957883875294,
3833=>456.55446984472434,
3834=>457.61384214488186,
3835=>458.6739027939789,
3836=>459.73464929637214,
3837=>460.7960791548032,
3838=>461.85818987040517,
3839=>462.9209789427081,
3840=>463.9844438696445,
3841=>465.0485821475575,
3842=>466.1133912712034,
3843=>467.1788687337594,
3844=>468.2450120268295,
3845=>469.3118186404501,
3846=>470.3792860630961,
3847=>471.4474117816866,
3848=>472.5161932815908,
3849=>473.5856280466342,
3850=>474.6557135591043,
3851=>475.7264472997566,
3852=>476.79782674782047,
3853=>477.8698493810044,
3854=>478.9425126755049,
3855=>480.01581410600784,
3856=>481.08975114569773,
3857=>482.1643212662627,
3858=>483.2395219379001,
3859=>484.31535062932335,
3860=>485.3918048077669,
3861=>486.4688819389928,
3862=>487.54657948729664,
3863=>488.6248949155132,
3864=>489.70382568502276,
3865=>490.7833692557569,
3866=>491.86352308620377,
3867=>492.9442846334169,
3868=>494.025651353017,
3869=>495.107620699201,
3870=>496.1901901247468,
3871=>497.2733570810196,
3872=>498.3571190179781,
3873=>499.4414733841799,
3874=>500.5264176267883,
3875=>501.61194919157754,
3876=>502.69806552293926,
3877=>503.7847640638885,
3878=>504.8720422560696,
3879=>505.95989753976227,
3880=>507.04832735388675,
3881=>508.137329136013,
3882=>509.2269003223622,
3883=>510.31703834781575,
3884=>511.40774064592057,
3885=>512.4990046488953,
3886=>513.5908277876358,
3887=>514.6832074917219,
3888=>515.7761411894231,
3889=>516.8696263077047,
3890=>517.9636602722337,
3891=>519.0582405073849,
3892=>520.1533644362473,
3893=>521.249029480629,
3894=>522.3452330610664,
3895=>523.4419725968261,
3896=>524.5392455059132,
3897=>525.6370492050773,
3898=>526.7353811098186,
3899=>527.8342386343936,
3900=>528.9336191918214,
3901=>530.0335201938898,
3902=>531.1339390511611,
3903=>532.2348731729786,
3904=>533.3363199674727,
3905=>534.4382768415667,
3906=>535.5407412009829,
3907=>536.6437104502493,
3908=>537.7471819927046,
3909=>538.8511532305056,
3910=>539.9556215646322,
3911=>541.0605843948946,
3912=>542.1660391199382,
3913=>543.2719831372508,
3914=>544.3784138431681,
3915=>545.4853286328799,
3916=>546.5927249004368,
3917=>547.7006000387546,
3918=>548.8089514396243,
3919=>549.9177764937132,
3920=>551.0270725905743,
3921=>552.136837118652,
3922=>553.2470674652873,
3923=>554.357761016725,
3924=>555.4689151581194,
3925=>556.5805272735402,
3926=>557.6925947459789,
3927=>558.8051149573552,
3928=>559.918085288523,
3929=>561.0315031192762,
3930=>562.1453658283554,
3931=>563.259670793453,
3932=>564.3744153912226,
3933=>565.4895969972802,
3934=>566.6052129862142,
3935=>567.7212607315901,
3936=>568.8377376059569,
3937=>569.9546409808536,
3938=>571.0719682268145,
3939=>572.1897167133769,
3940=>573.3078838090856,
3941=>574.4264668815002,
3942=>575.5454632972012,
3943=>576.6648704217955,
3944=>577.7846856199229,
3945=>578.9049062552642,
3946=>580.0255296905439,
3947=>581.1465532875386,
3948=>582.2679744070832,
3949=>583.3897904090763,
3950=>584.5119986524873,
3951=>585.6345964953617,
3952=>586.7575812948282,
3953=>587.8809504071044,
3954=>589.0047011875029,
3955=>590.128830990438,
3956=>591.2533371694317,
3957=>592.378217077119,
3958=>593.5034680652574,
3959=>594.6290874847284,
3960=>595.7550726855472,
3961=>596.8814210168676,
3962=>598.0081298269886,
3963=>599.1351964633603,
3964=>600.2626182725908,
3965=>601.3903926004517,
3966=>602.5185167918848,
3967=>603.6469881910085,
3968=>604.7758041411233,
3969=>605.9049619847187,
3970=>607.0344590634797,
3971=>608.1642927182913,
3972=>609.2944602892487,
3973=>610.4249591156588,
3974=>611.555786536049,
3975=>612.6869398881737,
3976=>613.8184165090195,
3977=>614.950213734812,
3978=>616.0823289010224,
3979=>617.2147593423729,
3980=>618.3475023928436,
3981=>619.4805553856789,
3982=>620.6139156533934,
3983=>621.7475805277779,
3984=>622.8815473399061,
3985=>624.0158134201424,
3986=>625.1503760981446,
3987=>626.2852327028734,
3988=>627.4203805625968,
3989=>628.5558170048978,
3990=>629.6915393566795,
3991=>630.8275449441724,
3992=>631.9638310929395,
3993=>633.100395127884,
3994=>634.2372343732544,
3995=>635.3743461526517,
3996=>636.5117277890347,
3997=>637.6493766047275,
3998=>638.7872899214244,
3999=>639.9254650601985,
4000=>641.0638993415051,
4001=>642.2025900851899,
4002=>643.3415346104946,
4003=>644.4807302360638,
4004=>645.6201742799506,
4005=>646.7598640596235,
4006=>647.8997968919725,
4007=>649.0399700933152,
4008=>650.1803809794035,
4009=>651.3210268654295,
4010=>652.4619050660324,
4011=>653.6030128953033,
4012=>654.7443476667953,
4013=>655.8859066935248,
4014=>657.027687287981,
4015=>658.1696867621317,
4016=>659.311902427429,
4017=>660.4543315948164,
4018=>661.5969715747344,
4019=>662.7398196771277,
4020=>663.8828732114505,
4021=>665.0261294866738,
4022=>666.1695858112909,
4023=>667.3132394933244,
4024=>668.4570878403323,
4025=>669.6011281594134,
4026=>670.7453577572169,
4027=>671.889773939944,
4028=>673.0343740133576,
4029=>674.1791552827875,
4030=>675.324115053137,
4031=>676.4692506288892,
4032=>677.614559314114,
4033=>678.7600384124714,
4034=>679.9056852272229,
4035=>681.051497061233,
4036=>682.1974712169804,
4037=>683.3436049965593,
4038=>684.4898957016887,
4039=>685.6363406337186,
4040=>686.7829370936354,
4041=>687.929682382069,
4042=>689.076573799299,
4043=>690.2236086452607,
4044=>691.3707842195522,
4045=>692.5180978214397,
4046=>693.6655467498649,
4047=>694.8131283034509,
4048=>695.9608397805081,
4049=>697.1086784790409,
4050=>698.2566416967561,
4051=>699.404726731065,
4052=>700.5529308790931,
4053=>701.7012514376853,
4054=>702.8496857034127,
4055=>703.9982309725784,
4056=>705.1468845412244,
4057=>706.2956437051376,
4058=>707.4445057598564,
4059=>708.5934680006767,
4060=>709.742527722659,
4061=>710.891682220634,
4062=>712.0409287892086,
4063=>713.190264722775,
4064=>714.3396873155132,
4065=>715.4891938613994,
4066=>716.6387816542126,
4067=>717.7884479875403,
4068=>718.9381901547852,
4069=>720.0880054491713,
4070=>721.2378911637506,
4071=>722.3878445914094,
4072=>723.5378630248742,
4073=>724.6879437567189,
4074=>725.8380840793706,
4075=>726.9882812851151,
4076=>728.1385326661069,
4077=>729.2888355143706,
4078=>730.43918712181,
4079=>731.5895847802149,
4080=>732.7400257812659,
4081=>733.8905074165419,
4082=>735.0410269775264,
4083=>736.191581755613,
4084=>737.3421690421129,
4085=>738.4927861282607,
4086=>739.6434303052205,
4087=>740.7940988640929,
4088=>741.9447890959212,
4089=>743.0954982916969,
4090=>744.2462237423687,
4091=>745.3969627388451,
4092=>746.5477125720035,
4093=>747.6984705326958,
4094=>748.8492339117546,
4095=>749.9999999999998
    );

signal lut_sig : unsigned(15 downto 0);

begin 
    sine <= STD_LOGIC_VECTOR(lut_sig);
    process (address)
            begin
                case address is
                   when x"000" => lut_sig <= to_unsigned(integer(my_rom(0)),16);
when x"001" => lut_sig <= to_unsigned(integer(my_rom(1)),16);
when x"002" => lut_sig <= to_unsigned(integer(my_rom(2)),16);
when x"003" => lut_sig <= to_unsigned(integer(my_rom(3)),16);
when x"004" => lut_sig <= to_unsigned(integer(my_rom(4)),16);
when x"005" => lut_sig <= to_unsigned(integer(my_rom(5)),16);
when x"006" => lut_sig <= to_unsigned(integer(my_rom(6)),16);
when x"007" => lut_sig <= to_unsigned(integer(my_rom(7)),16);
when x"008" => lut_sig <= to_unsigned(integer(my_rom(8)),16);
when x"009" => lut_sig <= to_unsigned(integer(my_rom(9)),16);
when x"00a" => lut_sig <= to_unsigned(integer(my_rom(10)),16);
when x"00b" => lut_sig <= to_unsigned(integer(my_rom(11)),16);
when x"00c" => lut_sig <= to_unsigned(integer(my_rom(12)),16);
when x"00d" => lut_sig <= to_unsigned(integer(my_rom(13)),16);
when x"00e" => lut_sig <= to_unsigned(integer(my_rom(14)),16);
when x"00f" => lut_sig <= to_unsigned(integer(my_rom(15)),16);
when x"010" => lut_sig <= to_unsigned(integer(my_rom(16)),16);
when x"011" => lut_sig <= to_unsigned(integer(my_rom(17)),16);
when x"012" => lut_sig <= to_unsigned(integer(my_rom(18)),16);
when x"013" => lut_sig <= to_unsigned(integer(my_rom(19)),16);
when x"014" => lut_sig <= to_unsigned(integer(my_rom(20)),16);
when x"015" => lut_sig <= to_unsigned(integer(my_rom(21)),16);
when x"016" => lut_sig <= to_unsigned(integer(my_rom(22)),16);
when x"017" => lut_sig <= to_unsigned(integer(my_rom(23)),16);
when x"018" => lut_sig <= to_unsigned(integer(my_rom(24)),16);
when x"019" => lut_sig <= to_unsigned(integer(my_rom(25)),16);
when x"01a" => lut_sig <= to_unsigned(integer(my_rom(26)),16);
when x"01b" => lut_sig <= to_unsigned(integer(my_rom(27)),16);
when x"01c" => lut_sig <= to_unsigned(integer(my_rom(28)),16);
when x"01d" => lut_sig <= to_unsigned(integer(my_rom(29)),16);
when x"01e" => lut_sig <= to_unsigned(integer(my_rom(30)),16);
when x"01f" => lut_sig <= to_unsigned(integer(my_rom(31)),16);
when x"020" => lut_sig <= to_unsigned(integer(my_rom(32)),16);
when x"021" => lut_sig <= to_unsigned(integer(my_rom(33)),16);
when x"022" => lut_sig <= to_unsigned(integer(my_rom(34)),16);
when x"023" => lut_sig <= to_unsigned(integer(my_rom(35)),16);
when x"024" => lut_sig <= to_unsigned(integer(my_rom(36)),16);
when x"025" => lut_sig <= to_unsigned(integer(my_rom(37)),16);
when x"026" => lut_sig <= to_unsigned(integer(my_rom(38)),16);
when x"027" => lut_sig <= to_unsigned(integer(my_rom(39)),16);
when x"028" => lut_sig <= to_unsigned(integer(my_rom(40)),16);
when x"029" => lut_sig <= to_unsigned(integer(my_rom(41)),16);
when x"02a" => lut_sig <= to_unsigned(integer(my_rom(42)),16);
when x"02b" => lut_sig <= to_unsigned(integer(my_rom(43)),16);
when x"02c" => lut_sig <= to_unsigned(integer(my_rom(44)),16);
when x"02d" => lut_sig <= to_unsigned(integer(my_rom(45)),16);
when x"02e" => lut_sig <= to_unsigned(integer(my_rom(46)),16);
when x"02f" => lut_sig <= to_unsigned(integer(my_rom(47)),16);
when x"030" => lut_sig <= to_unsigned(integer(my_rom(48)),16);
when x"031" => lut_sig <= to_unsigned(integer(my_rom(49)),16);
when x"032" => lut_sig <= to_unsigned(integer(my_rom(50)),16);
when x"033" => lut_sig <= to_unsigned(integer(my_rom(51)),16);
when x"034" => lut_sig <= to_unsigned(integer(my_rom(52)),16);
when x"035" => lut_sig <= to_unsigned(integer(my_rom(53)),16);
when x"036" => lut_sig <= to_unsigned(integer(my_rom(54)),16);
when x"037" => lut_sig <= to_unsigned(integer(my_rom(55)),16);
when x"038" => lut_sig <= to_unsigned(integer(my_rom(56)),16);
when x"039" => lut_sig <= to_unsigned(integer(my_rom(57)),16);
when x"03a" => lut_sig <= to_unsigned(integer(my_rom(58)),16);
when x"03b" => lut_sig <= to_unsigned(integer(my_rom(59)),16);
when x"03c" => lut_sig <= to_unsigned(integer(my_rom(60)),16);
when x"03d" => lut_sig <= to_unsigned(integer(my_rom(61)),16);
when x"03e" => lut_sig <= to_unsigned(integer(my_rom(62)),16);
when x"03f" => lut_sig <= to_unsigned(integer(my_rom(63)),16);
when x"040" => lut_sig <= to_unsigned(integer(my_rom(64)),16);
when x"041" => lut_sig <= to_unsigned(integer(my_rom(65)),16);
when x"042" => lut_sig <= to_unsigned(integer(my_rom(66)),16);
when x"043" => lut_sig <= to_unsigned(integer(my_rom(67)),16);
when x"044" => lut_sig <= to_unsigned(integer(my_rom(68)),16);
when x"045" => lut_sig <= to_unsigned(integer(my_rom(69)),16);
when x"046" => lut_sig <= to_unsigned(integer(my_rom(70)),16);
when x"047" => lut_sig <= to_unsigned(integer(my_rom(71)),16);
when x"048" => lut_sig <= to_unsigned(integer(my_rom(72)),16);
when x"049" => lut_sig <= to_unsigned(integer(my_rom(73)),16);
when x"04a" => lut_sig <= to_unsigned(integer(my_rom(74)),16);
when x"04b" => lut_sig <= to_unsigned(integer(my_rom(75)),16);
when x"04c" => lut_sig <= to_unsigned(integer(my_rom(76)),16);
when x"04d" => lut_sig <= to_unsigned(integer(my_rom(77)),16);
when x"04e" => lut_sig <= to_unsigned(integer(my_rom(78)),16);
when x"04f" => lut_sig <= to_unsigned(integer(my_rom(79)),16);
when x"050" => lut_sig <= to_unsigned(integer(my_rom(80)),16);
when x"051" => lut_sig <= to_unsigned(integer(my_rom(81)),16);
when x"052" => lut_sig <= to_unsigned(integer(my_rom(82)),16);
when x"053" => lut_sig <= to_unsigned(integer(my_rom(83)),16);
when x"054" => lut_sig <= to_unsigned(integer(my_rom(84)),16);
when x"055" => lut_sig <= to_unsigned(integer(my_rom(85)),16);
when x"056" => lut_sig <= to_unsigned(integer(my_rom(86)),16);
when x"057" => lut_sig <= to_unsigned(integer(my_rom(87)),16);
when x"058" => lut_sig <= to_unsigned(integer(my_rom(88)),16);
when x"059" => lut_sig <= to_unsigned(integer(my_rom(89)),16);
when x"05a" => lut_sig <= to_unsigned(integer(my_rom(90)),16);
when x"05b" => lut_sig <= to_unsigned(integer(my_rom(91)),16);
when x"05c" => lut_sig <= to_unsigned(integer(my_rom(92)),16);
when x"05d" => lut_sig <= to_unsigned(integer(my_rom(93)),16);
when x"05e" => lut_sig <= to_unsigned(integer(my_rom(94)),16);
when x"05f" => lut_sig <= to_unsigned(integer(my_rom(95)),16);
when x"060" => lut_sig <= to_unsigned(integer(my_rom(96)),16);
when x"061" => lut_sig <= to_unsigned(integer(my_rom(97)),16);
when x"062" => lut_sig <= to_unsigned(integer(my_rom(98)),16);
when x"063" => lut_sig <= to_unsigned(integer(my_rom(99)),16);
when x"064" => lut_sig <= to_unsigned(integer(my_rom(100)),16);
when x"065" => lut_sig <= to_unsigned(integer(my_rom(101)),16);
when x"066" => lut_sig <= to_unsigned(integer(my_rom(102)),16);
when x"067" => lut_sig <= to_unsigned(integer(my_rom(103)),16);
when x"068" => lut_sig <= to_unsigned(integer(my_rom(104)),16);
when x"069" => lut_sig <= to_unsigned(integer(my_rom(105)),16);
when x"06a" => lut_sig <= to_unsigned(integer(my_rom(106)),16);
when x"06b" => lut_sig <= to_unsigned(integer(my_rom(107)),16);
when x"06c" => lut_sig <= to_unsigned(integer(my_rom(108)),16);
when x"06d" => lut_sig <= to_unsigned(integer(my_rom(109)),16);
when x"06e" => lut_sig <= to_unsigned(integer(my_rom(110)),16);
when x"06f" => lut_sig <= to_unsigned(integer(my_rom(111)),16);
when x"070" => lut_sig <= to_unsigned(integer(my_rom(112)),16);
when x"071" => lut_sig <= to_unsigned(integer(my_rom(113)),16);
when x"072" => lut_sig <= to_unsigned(integer(my_rom(114)),16);
when x"073" => lut_sig <= to_unsigned(integer(my_rom(115)),16);
when x"074" => lut_sig <= to_unsigned(integer(my_rom(116)),16);
when x"075" => lut_sig <= to_unsigned(integer(my_rom(117)),16);
when x"076" => lut_sig <= to_unsigned(integer(my_rom(118)),16);
when x"077" => lut_sig <= to_unsigned(integer(my_rom(119)),16);
when x"078" => lut_sig <= to_unsigned(integer(my_rom(120)),16);
when x"079" => lut_sig <= to_unsigned(integer(my_rom(121)),16);
when x"07a" => lut_sig <= to_unsigned(integer(my_rom(122)),16);
when x"07b" => lut_sig <= to_unsigned(integer(my_rom(123)),16);
when x"07c" => lut_sig <= to_unsigned(integer(my_rom(124)),16);
when x"07d" => lut_sig <= to_unsigned(integer(my_rom(125)),16);
when x"07e" => lut_sig <= to_unsigned(integer(my_rom(126)),16);
when x"07f" => lut_sig <= to_unsigned(integer(my_rom(127)),16);
when x"080" => lut_sig <= to_unsigned(integer(my_rom(128)),16);
when x"081" => lut_sig <= to_unsigned(integer(my_rom(129)),16);
when x"082" => lut_sig <= to_unsigned(integer(my_rom(130)),16);
when x"083" => lut_sig <= to_unsigned(integer(my_rom(131)),16);
when x"084" => lut_sig <= to_unsigned(integer(my_rom(132)),16);
when x"085" => lut_sig <= to_unsigned(integer(my_rom(133)),16);
when x"086" => lut_sig <= to_unsigned(integer(my_rom(134)),16);
when x"087" => lut_sig <= to_unsigned(integer(my_rom(135)),16);
when x"088" => lut_sig <= to_unsigned(integer(my_rom(136)),16);
when x"089" => lut_sig <= to_unsigned(integer(my_rom(137)),16);
when x"08a" => lut_sig <= to_unsigned(integer(my_rom(138)),16);
when x"08b" => lut_sig <= to_unsigned(integer(my_rom(139)),16);
when x"08c" => lut_sig <= to_unsigned(integer(my_rom(140)),16);
when x"08d" => lut_sig <= to_unsigned(integer(my_rom(141)),16);
when x"08e" => lut_sig <= to_unsigned(integer(my_rom(142)),16);
when x"08f" => lut_sig <= to_unsigned(integer(my_rom(143)),16);
when x"090" => lut_sig <= to_unsigned(integer(my_rom(144)),16);
when x"091" => lut_sig <= to_unsigned(integer(my_rom(145)),16);
when x"092" => lut_sig <= to_unsigned(integer(my_rom(146)),16);
when x"093" => lut_sig <= to_unsigned(integer(my_rom(147)),16);
when x"094" => lut_sig <= to_unsigned(integer(my_rom(148)),16);
when x"095" => lut_sig <= to_unsigned(integer(my_rom(149)),16);
when x"096" => lut_sig <= to_unsigned(integer(my_rom(150)),16);
when x"097" => lut_sig <= to_unsigned(integer(my_rom(151)),16);
when x"098" => lut_sig <= to_unsigned(integer(my_rom(152)),16);
when x"099" => lut_sig <= to_unsigned(integer(my_rom(153)),16);
when x"09a" => lut_sig <= to_unsigned(integer(my_rom(154)),16);
when x"09b" => lut_sig <= to_unsigned(integer(my_rom(155)),16);
when x"09c" => lut_sig <= to_unsigned(integer(my_rom(156)),16);
when x"09d" => lut_sig <= to_unsigned(integer(my_rom(157)),16);
when x"09e" => lut_sig <= to_unsigned(integer(my_rom(158)),16);
when x"09f" => lut_sig <= to_unsigned(integer(my_rom(159)),16);
when x"0a0" => lut_sig <= to_unsigned(integer(my_rom(160)),16);
when x"0a1" => lut_sig <= to_unsigned(integer(my_rom(161)),16);
when x"0a2" => lut_sig <= to_unsigned(integer(my_rom(162)),16);
when x"0a3" => lut_sig <= to_unsigned(integer(my_rom(163)),16);
when x"0a4" => lut_sig <= to_unsigned(integer(my_rom(164)),16);
when x"0a5" => lut_sig <= to_unsigned(integer(my_rom(165)),16);
when x"0a6" => lut_sig <= to_unsigned(integer(my_rom(166)),16);
when x"0a7" => lut_sig <= to_unsigned(integer(my_rom(167)),16);
when x"0a8" => lut_sig <= to_unsigned(integer(my_rom(168)),16);
when x"0a9" => lut_sig <= to_unsigned(integer(my_rom(169)),16);
when x"0aa" => lut_sig <= to_unsigned(integer(my_rom(170)),16);
when x"0ab" => lut_sig <= to_unsigned(integer(my_rom(171)),16);
when x"0ac" => lut_sig <= to_unsigned(integer(my_rom(172)),16);
when x"0ad" => lut_sig <= to_unsigned(integer(my_rom(173)),16);
when x"0ae" => lut_sig <= to_unsigned(integer(my_rom(174)),16);
when x"0af" => lut_sig <= to_unsigned(integer(my_rom(175)),16);
when x"0b0" => lut_sig <= to_unsigned(integer(my_rom(176)),16);
when x"0b1" => lut_sig <= to_unsigned(integer(my_rom(177)),16);
when x"0b2" => lut_sig <= to_unsigned(integer(my_rom(178)),16);
when x"0b3" => lut_sig <= to_unsigned(integer(my_rom(179)),16);
when x"0b4" => lut_sig <= to_unsigned(integer(my_rom(180)),16);
when x"0b5" => lut_sig <= to_unsigned(integer(my_rom(181)),16);
when x"0b6" => lut_sig <= to_unsigned(integer(my_rom(182)),16);
when x"0b7" => lut_sig <= to_unsigned(integer(my_rom(183)),16);
when x"0b8" => lut_sig <= to_unsigned(integer(my_rom(184)),16);
when x"0b9" => lut_sig <= to_unsigned(integer(my_rom(185)),16);
when x"0ba" => lut_sig <= to_unsigned(integer(my_rom(186)),16);
when x"0bb" => lut_sig <= to_unsigned(integer(my_rom(187)),16);
when x"0bc" => lut_sig <= to_unsigned(integer(my_rom(188)),16);
when x"0bd" => lut_sig <= to_unsigned(integer(my_rom(189)),16);
when x"0be" => lut_sig <= to_unsigned(integer(my_rom(190)),16);
when x"0bf" => lut_sig <= to_unsigned(integer(my_rom(191)),16);
when x"0c0" => lut_sig <= to_unsigned(integer(my_rom(192)),16);
when x"0c1" => lut_sig <= to_unsigned(integer(my_rom(193)),16);
when x"0c2" => lut_sig <= to_unsigned(integer(my_rom(194)),16);
when x"0c3" => lut_sig <= to_unsigned(integer(my_rom(195)),16);
when x"0c4" => lut_sig <= to_unsigned(integer(my_rom(196)),16);
when x"0c5" => lut_sig <= to_unsigned(integer(my_rom(197)),16);
when x"0c6" => lut_sig <= to_unsigned(integer(my_rom(198)),16);
when x"0c7" => lut_sig <= to_unsigned(integer(my_rom(199)),16);
when x"0c8" => lut_sig <= to_unsigned(integer(my_rom(200)),16);
when x"0c9" => lut_sig <= to_unsigned(integer(my_rom(201)),16);
when x"0ca" => lut_sig <= to_unsigned(integer(my_rom(202)),16);
when x"0cb" => lut_sig <= to_unsigned(integer(my_rom(203)),16);
when x"0cc" => lut_sig <= to_unsigned(integer(my_rom(204)),16);
when x"0cd" => lut_sig <= to_unsigned(integer(my_rom(205)),16);
when x"0ce" => lut_sig <= to_unsigned(integer(my_rom(206)),16);
when x"0cf" => lut_sig <= to_unsigned(integer(my_rom(207)),16);
when x"0d0" => lut_sig <= to_unsigned(integer(my_rom(208)),16);
when x"0d1" => lut_sig <= to_unsigned(integer(my_rom(209)),16);
when x"0d2" => lut_sig <= to_unsigned(integer(my_rom(210)),16);
when x"0d3" => lut_sig <= to_unsigned(integer(my_rom(211)),16);
when x"0d4" => lut_sig <= to_unsigned(integer(my_rom(212)),16);
when x"0d5" => lut_sig <= to_unsigned(integer(my_rom(213)),16);
when x"0d6" => lut_sig <= to_unsigned(integer(my_rom(214)),16);
when x"0d7" => lut_sig <= to_unsigned(integer(my_rom(215)),16);
when x"0d8" => lut_sig <= to_unsigned(integer(my_rom(216)),16);
when x"0d9" => lut_sig <= to_unsigned(integer(my_rom(217)),16);
when x"0da" => lut_sig <= to_unsigned(integer(my_rom(218)),16);
when x"0db" => lut_sig <= to_unsigned(integer(my_rom(219)),16);
when x"0dc" => lut_sig <= to_unsigned(integer(my_rom(220)),16);
when x"0dd" => lut_sig <= to_unsigned(integer(my_rom(221)),16);
when x"0de" => lut_sig <= to_unsigned(integer(my_rom(222)),16);
when x"0df" => lut_sig <= to_unsigned(integer(my_rom(223)),16);
when x"0e0" => lut_sig <= to_unsigned(integer(my_rom(224)),16);
when x"0e1" => lut_sig <= to_unsigned(integer(my_rom(225)),16);
when x"0e2" => lut_sig <= to_unsigned(integer(my_rom(226)),16);
when x"0e3" => lut_sig <= to_unsigned(integer(my_rom(227)),16);
when x"0e4" => lut_sig <= to_unsigned(integer(my_rom(228)),16);
when x"0e5" => lut_sig <= to_unsigned(integer(my_rom(229)),16);
when x"0e6" => lut_sig <= to_unsigned(integer(my_rom(230)),16);
when x"0e7" => lut_sig <= to_unsigned(integer(my_rom(231)),16);
when x"0e8" => lut_sig <= to_unsigned(integer(my_rom(232)),16);
when x"0e9" => lut_sig <= to_unsigned(integer(my_rom(233)),16);
when x"0ea" => lut_sig <= to_unsigned(integer(my_rom(234)),16);
when x"0eb" => lut_sig <= to_unsigned(integer(my_rom(235)),16);
when x"0ec" => lut_sig <= to_unsigned(integer(my_rom(236)),16);
when x"0ed" => lut_sig <= to_unsigned(integer(my_rom(237)),16);
when x"0ee" => lut_sig <= to_unsigned(integer(my_rom(238)),16);
when x"0ef" => lut_sig <= to_unsigned(integer(my_rom(239)),16);
when x"0f0" => lut_sig <= to_unsigned(integer(my_rom(240)),16);
when x"0f1" => lut_sig <= to_unsigned(integer(my_rom(241)),16);
when x"0f2" => lut_sig <= to_unsigned(integer(my_rom(242)),16);
when x"0f3" => lut_sig <= to_unsigned(integer(my_rom(243)),16);
when x"0f4" => lut_sig <= to_unsigned(integer(my_rom(244)),16);
when x"0f5" => lut_sig <= to_unsigned(integer(my_rom(245)),16);
when x"0f6" => lut_sig <= to_unsigned(integer(my_rom(246)),16);
when x"0f7" => lut_sig <= to_unsigned(integer(my_rom(247)),16);
when x"0f8" => lut_sig <= to_unsigned(integer(my_rom(248)),16);
when x"0f9" => lut_sig <= to_unsigned(integer(my_rom(249)),16);
when x"0fa" => lut_sig <= to_unsigned(integer(my_rom(250)),16);
when x"0fb" => lut_sig <= to_unsigned(integer(my_rom(251)),16);
when x"0fc" => lut_sig <= to_unsigned(integer(my_rom(252)),16);
when x"0fd" => lut_sig <= to_unsigned(integer(my_rom(253)),16);
when x"0fe" => lut_sig <= to_unsigned(integer(my_rom(254)),16);
when x"0ff" => lut_sig <= to_unsigned(integer(my_rom(255)),16);
when x"100" => lut_sig <= to_unsigned(integer(my_rom(256)),16);
when x"101" => lut_sig <= to_unsigned(integer(my_rom(257)),16);
when x"102" => lut_sig <= to_unsigned(integer(my_rom(258)),16);
when x"103" => lut_sig <= to_unsigned(integer(my_rom(259)),16);
when x"104" => lut_sig <= to_unsigned(integer(my_rom(260)),16);
when x"105" => lut_sig <= to_unsigned(integer(my_rom(261)),16);
when x"106" => lut_sig <= to_unsigned(integer(my_rom(262)),16);
when x"107" => lut_sig <= to_unsigned(integer(my_rom(263)),16);
when x"108" => lut_sig <= to_unsigned(integer(my_rom(264)),16);
when x"109" => lut_sig <= to_unsigned(integer(my_rom(265)),16);
when x"10a" => lut_sig <= to_unsigned(integer(my_rom(266)),16);
when x"10b" => lut_sig <= to_unsigned(integer(my_rom(267)),16);
when x"10c" => lut_sig <= to_unsigned(integer(my_rom(268)),16);
when x"10d" => lut_sig <= to_unsigned(integer(my_rom(269)),16);
when x"10e" => lut_sig <= to_unsigned(integer(my_rom(270)),16);
when x"10f" => lut_sig <= to_unsigned(integer(my_rom(271)),16);
when x"110" => lut_sig <= to_unsigned(integer(my_rom(272)),16);
when x"111" => lut_sig <= to_unsigned(integer(my_rom(273)),16);
when x"112" => lut_sig <= to_unsigned(integer(my_rom(274)),16);
when x"113" => lut_sig <= to_unsigned(integer(my_rom(275)),16);
when x"114" => lut_sig <= to_unsigned(integer(my_rom(276)),16);
when x"115" => lut_sig <= to_unsigned(integer(my_rom(277)),16);
when x"116" => lut_sig <= to_unsigned(integer(my_rom(278)),16);
when x"117" => lut_sig <= to_unsigned(integer(my_rom(279)),16);
when x"118" => lut_sig <= to_unsigned(integer(my_rom(280)),16);
when x"119" => lut_sig <= to_unsigned(integer(my_rom(281)),16);
when x"11a" => lut_sig <= to_unsigned(integer(my_rom(282)),16);
when x"11b" => lut_sig <= to_unsigned(integer(my_rom(283)),16);
when x"11c" => lut_sig <= to_unsigned(integer(my_rom(284)),16);
when x"11d" => lut_sig <= to_unsigned(integer(my_rom(285)),16);
when x"11e" => lut_sig <= to_unsigned(integer(my_rom(286)),16);
when x"11f" => lut_sig <= to_unsigned(integer(my_rom(287)),16);
when x"120" => lut_sig <= to_unsigned(integer(my_rom(288)),16);
when x"121" => lut_sig <= to_unsigned(integer(my_rom(289)),16);
when x"122" => lut_sig <= to_unsigned(integer(my_rom(290)),16);
when x"123" => lut_sig <= to_unsigned(integer(my_rom(291)),16);
when x"124" => lut_sig <= to_unsigned(integer(my_rom(292)),16);
when x"125" => lut_sig <= to_unsigned(integer(my_rom(293)),16);
when x"126" => lut_sig <= to_unsigned(integer(my_rom(294)),16);
when x"127" => lut_sig <= to_unsigned(integer(my_rom(295)),16);
when x"128" => lut_sig <= to_unsigned(integer(my_rom(296)),16);
when x"129" => lut_sig <= to_unsigned(integer(my_rom(297)),16);
when x"12a" => lut_sig <= to_unsigned(integer(my_rom(298)),16);
when x"12b" => lut_sig <= to_unsigned(integer(my_rom(299)),16);
when x"12c" => lut_sig <= to_unsigned(integer(my_rom(300)),16);
when x"12d" => lut_sig <= to_unsigned(integer(my_rom(301)),16);
when x"12e" => lut_sig <= to_unsigned(integer(my_rom(302)),16);
when x"12f" => lut_sig <= to_unsigned(integer(my_rom(303)),16);
when x"130" => lut_sig <= to_unsigned(integer(my_rom(304)),16);
when x"131" => lut_sig <= to_unsigned(integer(my_rom(305)),16);
when x"132" => lut_sig <= to_unsigned(integer(my_rom(306)),16);
when x"133" => lut_sig <= to_unsigned(integer(my_rom(307)),16);
when x"134" => lut_sig <= to_unsigned(integer(my_rom(308)),16);
when x"135" => lut_sig <= to_unsigned(integer(my_rom(309)),16);
when x"136" => lut_sig <= to_unsigned(integer(my_rom(310)),16);
when x"137" => lut_sig <= to_unsigned(integer(my_rom(311)),16);
when x"138" => lut_sig <= to_unsigned(integer(my_rom(312)),16);
when x"139" => lut_sig <= to_unsigned(integer(my_rom(313)),16);
when x"13a" => lut_sig <= to_unsigned(integer(my_rom(314)),16);
when x"13b" => lut_sig <= to_unsigned(integer(my_rom(315)),16);
when x"13c" => lut_sig <= to_unsigned(integer(my_rom(316)),16);
when x"13d" => lut_sig <= to_unsigned(integer(my_rom(317)),16);
when x"13e" => lut_sig <= to_unsigned(integer(my_rom(318)),16);
when x"13f" => lut_sig <= to_unsigned(integer(my_rom(319)),16);
when x"140" => lut_sig <= to_unsigned(integer(my_rom(320)),16);
when x"141" => lut_sig <= to_unsigned(integer(my_rom(321)),16);
when x"142" => lut_sig <= to_unsigned(integer(my_rom(322)),16);
when x"143" => lut_sig <= to_unsigned(integer(my_rom(323)),16);
when x"144" => lut_sig <= to_unsigned(integer(my_rom(324)),16);
when x"145" => lut_sig <= to_unsigned(integer(my_rom(325)),16);
when x"146" => lut_sig <= to_unsigned(integer(my_rom(326)),16);
when x"147" => lut_sig <= to_unsigned(integer(my_rom(327)),16);
when x"148" => lut_sig <= to_unsigned(integer(my_rom(328)),16);
when x"149" => lut_sig <= to_unsigned(integer(my_rom(329)),16);
when x"14a" => lut_sig <= to_unsigned(integer(my_rom(330)),16);
when x"14b" => lut_sig <= to_unsigned(integer(my_rom(331)),16);
when x"14c" => lut_sig <= to_unsigned(integer(my_rom(332)),16);
when x"14d" => lut_sig <= to_unsigned(integer(my_rom(333)),16);
when x"14e" => lut_sig <= to_unsigned(integer(my_rom(334)),16);
when x"14f" => lut_sig <= to_unsigned(integer(my_rom(335)),16);
when x"150" => lut_sig <= to_unsigned(integer(my_rom(336)),16);
when x"151" => lut_sig <= to_unsigned(integer(my_rom(337)),16);
when x"152" => lut_sig <= to_unsigned(integer(my_rom(338)),16);
when x"153" => lut_sig <= to_unsigned(integer(my_rom(339)),16);
when x"154" => lut_sig <= to_unsigned(integer(my_rom(340)),16);
when x"155" => lut_sig <= to_unsigned(integer(my_rom(341)),16);
when x"156" => lut_sig <= to_unsigned(integer(my_rom(342)),16);
when x"157" => lut_sig <= to_unsigned(integer(my_rom(343)),16);
when x"158" => lut_sig <= to_unsigned(integer(my_rom(344)),16);
when x"159" => lut_sig <= to_unsigned(integer(my_rom(345)),16);
when x"15a" => lut_sig <= to_unsigned(integer(my_rom(346)),16);
when x"15b" => lut_sig <= to_unsigned(integer(my_rom(347)),16);
when x"15c" => lut_sig <= to_unsigned(integer(my_rom(348)),16);
when x"15d" => lut_sig <= to_unsigned(integer(my_rom(349)),16);
when x"15e" => lut_sig <= to_unsigned(integer(my_rom(350)),16);
when x"15f" => lut_sig <= to_unsigned(integer(my_rom(351)),16);
when x"160" => lut_sig <= to_unsigned(integer(my_rom(352)),16);
when x"161" => lut_sig <= to_unsigned(integer(my_rom(353)),16);
when x"162" => lut_sig <= to_unsigned(integer(my_rom(354)),16);
when x"163" => lut_sig <= to_unsigned(integer(my_rom(355)),16);
when x"164" => lut_sig <= to_unsigned(integer(my_rom(356)),16);
when x"165" => lut_sig <= to_unsigned(integer(my_rom(357)),16);
when x"166" => lut_sig <= to_unsigned(integer(my_rom(358)),16);
when x"167" => lut_sig <= to_unsigned(integer(my_rom(359)),16);
when x"168" => lut_sig <= to_unsigned(integer(my_rom(360)),16);
when x"169" => lut_sig <= to_unsigned(integer(my_rom(361)),16);
when x"16a" => lut_sig <= to_unsigned(integer(my_rom(362)),16);
when x"16b" => lut_sig <= to_unsigned(integer(my_rom(363)),16);
when x"16c" => lut_sig <= to_unsigned(integer(my_rom(364)),16);
when x"16d" => lut_sig <= to_unsigned(integer(my_rom(365)),16);
when x"16e" => lut_sig <= to_unsigned(integer(my_rom(366)),16);
when x"16f" => lut_sig <= to_unsigned(integer(my_rom(367)),16);
when x"170" => lut_sig <= to_unsigned(integer(my_rom(368)),16);
when x"171" => lut_sig <= to_unsigned(integer(my_rom(369)),16);
when x"172" => lut_sig <= to_unsigned(integer(my_rom(370)),16);
when x"173" => lut_sig <= to_unsigned(integer(my_rom(371)),16);
when x"174" => lut_sig <= to_unsigned(integer(my_rom(372)),16);
when x"175" => lut_sig <= to_unsigned(integer(my_rom(373)),16);
when x"176" => lut_sig <= to_unsigned(integer(my_rom(374)),16);
when x"177" => lut_sig <= to_unsigned(integer(my_rom(375)),16);
when x"178" => lut_sig <= to_unsigned(integer(my_rom(376)),16);
when x"179" => lut_sig <= to_unsigned(integer(my_rom(377)),16);
when x"17a" => lut_sig <= to_unsigned(integer(my_rom(378)),16);
when x"17b" => lut_sig <= to_unsigned(integer(my_rom(379)),16);
when x"17c" => lut_sig <= to_unsigned(integer(my_rom(380)),16);
when x"17d" => lut_sig <= to_unsigned(integer(my_rom(381)),16);
when x"17e" => lut_sig <= to_unsigned(integer(my_rom(382)),16);
when x"17f" => lut_sig <= to_unsigned(integer(my_rom(383)),16);
when x"180" => lut_sig <= to_unsigned(integer(my_rom(384)),16);
when x"181" => lut_sig <= to_unsigned(integer(my_rom(385)),16);
when x"182" => lut_sig <= to_unsigned(integer(my_rom(386)),16);
when x"183" => lut_sig <= to_unsigned(integer(my_rom(387)),16);
when x"184" => lut_sig <= to_unsigned(integer(my_rom(388)),16);
when x"185" => lut_sig <= to_unsigned(integer(my_rom(389)),16);
when x"186" => lut_sig <= to_unsigned(integer(my_rom(390)),16);
when x"187" => lut_sig <= to_unsigned(integer(my_rom(391)),16);
when x"188" => lut_sig <= to_unsigned(integer(my_rom(392)),16);
when x"189" => lut_sig <= to_unsigned(integer(my_rom(393)),16);
when x"18a" => lut_sig <= to_unsigned(integer(my_rom(394)),16);
when x"18b" => lut_sig <= to_unsigned(integer(my_rom(395)),16);
when x"18c" => lut_sig <= to_unsigned(integer(my_rom(396)),16);
when x"18d" => lut_sig <= to_unsigned(integer(my_rom(397)),16);
when x"18e" => lut_sig <= to_unsigned(integer(my_rom(398)),16);
when x"18f" => lut_sig <= to_unsigned(integer(my_rom(399)),16);
when x"190" => lut_sig <= to_unsigned(integer(my_rom(400)),16);
when x"191" => lut_sig <= to_unsigned(integer(my_rom(401)),16);
when x"192" => lut_sig <= to_unsigned(integer(my_rom(402)),16);
when x"193" => lut_sig <= to_unsigned(integer(my_rom(403)),16);
when x"194" => lut_sig <= to_unsigned(integer(my_rom(404)),16);
when x"195" => lut_sig <= to_unsigned(integer(my_rom(405)),16);
when x"196" => lut_sig <= to_unsigned(integer(my_rom(406)),16);
when x"197" => lut_sig <= to_unsigned(integer(my_rom(407)),16);
when x"198" => lut_sig <= to_unsigned(integer(my_rom(408)),16);
when x"199" => lut_sig <= to_unsigned(integer(my_rom(409)),16);
when x"19a" => lut_sig <= to_unsigned(integer(my_rom(410)),16);
when x"19b" => lut_sig <= to_unsigned(integer(my_rom(411)),16);
when x"19c" => lut_sig <= to_unsigned(integer(my_rom(412)),16);
when x"19d" => lut_sig <= to_unsigned(integer(my_rom(413)),16);
when x"19e" => lut_sig <= to_unsigned(integer(my_rom(414)),16);
when x"19f" => lut_sig <= to_unsigned(integer(my_rom(415)),16);
when x"1a0" => lut_sig <= to_unsigned(integer(my_rom(416)),16);
when x"1a1" => lut_sig <= to_unsigned(integer(my_rom(417)),16);
when x"1a2" => lut_sig <= to_unsigned(integer(my_rom(418)),16);
when x"1a3" => lut_sig <= to_unsigned(integer(my_rom(419)),16);
when x"1a4" => lut_sig <= to_unsigned(integer(my_rom(420)),16);
when x"1a5" => lut_sig <= to_unsigned(integer(my_rom(421)),16);
when x"1a6" => lut_sig <= to_unsigned(integer(my_rom(422)),16);
when x"1a7" => lut_sig <= to_unsigned(integer(my_rom(423)),16);
when x"1a8" => lut_sig <= to_unsigned(integer(my_rom(424)),16);
when x"1a9" => lut_sig <= to_unsigned(integer(my_rom(425)),16);
when x"1aa" => lut_sig <= to_unsigned(integer(my_rom(426)),16);
when x"1ab" => lut_sig <= to_unsigned(integer(my_rom(427)),16);
when x"1ac" => lut_sig <= to_unsigned(integer(my_rom(428)),16);
when x"1ad" => lut_sig <= to_unsigned(integer(my_rom(429)),16);
when x"1ae" => lut_sig <= to_unsigned(integer(my_rom(430)),16);
when x"1af" => lut_sig <= to_unsigned(integer(my_rom(431)),16);
when x"1b0" => lut_sig <= to_unsigned(integer(my_rom(432)),16);
when x"1b1" => lut_sig <= to_unsigned(integer(my_rom(433)),16);
when x"1b2" => lut_sig <= to_unsigned(integer(my_rom(434)),16);
when x"1b3" => lut_sig <= to_unsigned(integer(my_rom(435)),16);
when x"1b4" => lut_sig <= to_unsigned(integer(my_rom(436)),16);
when x"1b5" => lut_sig <= to_unsigned(integer(my_rom(437)),16);
when x"1b6" => lut_sig <= to_unsigned(integer(my_rom(438)),16);
when x"1b7" => lut_sig <= to_unsigned(integer(my_rom(439)),16);
when x"1b8" => lut_sig <= to_unsigned(integer(my_rom(440)),16);
when x"1b9" => lut_sig <= to_unsigned(integer(my_rom(441)),16);
when x"1ba" => lut_sig <= to_unsigned(integer(my_rom(442)),16);
when x"1bb" => lut_sig <= to_unsigned(integer(my_rom(443)),16);
when x"1bc" => lut_sig <= to_unsigned(integer(my_rom(444)),16);
when x"1bd" => lut_sig <= to_unsigned(integer(my_rom(445)),16);
when x"1be" => lut_sig <= to_unsigned(integer(my_rom(446)),16);
when x"1bf" => lut_sig <= to_unsigned(integer(my_rom(447)),16);
when x"1c0" => lut_sig <= to_unsigned(integer(my_rom(448)),16);
when x"1c1" => lut_sig <= to_unsigned(integer(my_rom(449)),16);
when x"1c2" => lut_sig <= to_unsigned(integer(my_rom(450)),16);
when x"1c3" => lut_sig <= to_unsigned(integer(my_rom(451)),16);
when x"1c4" => lut_sig <= to_unsigned(integer(my_rom(452)),16);
when x"1c5" => lut_sig <= to_unsigned(integer(my_rom(453)),16);
when x"1c6" => lut_sig <= to_unsigned(integer(my_rom(454)),16);
when x"1c7" => lut_sig <= to_unsigned(integer(my_rom(455)),16);
when x"1c8" => lut_sig <= to_unsigned(integer(my_rom(456)),16);
when x"1c9" => lut_sig <= to_unsigned(integer(my_rom(457)),16);
when x"1ca" => lut_sig <= to_unsigned(integer(my_rom(458)),16);
when x"1cb" => lut_sig <= to_unsigned(integer(my_rom(459)),16);
when x"1cc" => lut_sig <= to_unsigned(integer(my_rom(460)),16);
when x"1cd" => lut_sig <= to_unsigned(integer(my_rom(461)),16);
when x"1ce" => lut_sig <= to_unsigned(integer(my_rom(462)),16);
when x"1cf" => lut_sig <= to_unsigned(integer(my_rom(463)),16);
when x"1d0" => lut_sig <= to_unsigned(integer(my_rom(464)),16);
when x"1d1" => lut_sig <= to_unsigned(integer(my_rom(465)),16);
when x"1d2" => lut_sig <= to_unsigned(integer(my_rom(466)),16);
when x"1d3" => lut_sig <= to_unsigned(integer(my_rom(467)),16);
when x"1d4" => lut_sig <= to_unsigned(integer(my_rom(468)),16);
when x"1d5" => lut_sig <= to_unsigned(integer(my_rom(469)),16);
when x"1d6" => lut_sig <= to_unsigned(integer(my_rom(470)),16);
when x"1d7" => lut_sig <= to_unsigned(integer(my_rom(471)),16);
when x"1d8" => lut_sig <= to_unsigned(integer(my_rom(472)),16);
when x"1d9" => lut_sig <= to_unsigned(integer(my_rom(473)),16);
when x"1da" => lut_sig <= to_unsigned(integer(my_rom(474)),16);
when x"1db" => lut_sig <= to_unsigned(integer(my_rom(475)),16);
when x"1dc" => lut_sig <= to_unsigned(integer(my_rom(476)),16);
when x"1dd" => lut_sig <= to_unsigned(integer(my_rom(477)),16);
when x"1de" => lut_sig <= to_unsigned(integer(my_rom(478)),16);
when x"1df" => lut_sig <= to_unsigned(integer(my_rom(479)),16);
when x"1e0" => lut_sig <= to_unsigned(integer(my_rom(480)),16);
when x"1e1" => lut_sig <= to_unsigned(integer(my_rom(481)),16);
when x"1e2" => lut_sig <= to_unsigned(integer(my_rom(482)),16);
when x"1e3" => lut_sig <= to_unsigned(integer(my_rom(483)),16);
when x"1e4" => lut_sig <= to_unsigned(integer(my_rom(484)),16);
when x"1e5" => lut_sig <= to_unsigned(integer(my_rom(485)),16);
when x"1e6" => lut_sig <= to_unsigned(integer(my_rom(486)),16);
when x"1e7" => lut_sig <= to_unsigned(integer(my_rom(487)),16);
when x"1e8" => lut_sig <= to_unsigned(integer(my_rom(488)),16);
when x"1e9" => lut_sig <= to_unsigned(integer(my_rom(489)),16);
when x"1ea" => lut_sig <= to_unsigned(integer(my_rom(490)),16);
when x"1eb" => lut_sig <= to_unsigned(integer(my_rom(491)),16);
when x"1ec" => lut_sig <= to_unsigned(integer(my_rom(492)),16);
when x"1ed" => lut_sig <= to_unsigned(integer(my_rom(493)),16);
when x"1ee" => lut_sig <= to_unsigned(integer(my_rom(494)),16);
when x"1ef" => lut_sig <= to_unsigned(integer(my_rom(495)),16);
when x"1f0" => lut_sig <= to_unsigned(integer(my_rom(496)),16);
when x"1f1" => lut_sig <= to_unsigned(integer(my_rom(497)),16);
when x"1f2" => lut_sig <= to_unsigned(integer(my_rom(498)),16);
when x"1f3" => lut_sig <= to_unsigned(integer(my_rom(499)),16);
when x"1f4" => lut_sig <= to_unsigned(integer(my_rom(500)),16);
when x"1f5" => lut_sig <= to_unsigned(integer(my_rom(501)),16);
when x"1f6" => lut_sig <= to_unsigned(integer(my_rom(502)),16);
when x"1f7" => lut_sig <= to_unsigned(integer(my_rom(503)),16);
when x"1f8" => lut_sig <= to_unsigned(integer(my_rom(504)),16);
when x"1f9" => lut_sig <= to_unsigned(integer(my_rom(505)),16);
when x"1fa" => lut_sig <= to_unsigned(integer(my_rom(506)),16);
when x"1fb" => lut_sig <= to_unsigned(integer(my_rom(507)),16);
when x"1fc" => lut_sig <= to_unsigned(integer(my_rom(508)),16);
when x"1fd" => lut_sig <= to_unsigned(integer(my_rom(509)),16);
when x"1fe" => lut_sig <= to_unsigned(integer(my_rom(510)),16);
when x"1ff" => lut_sig <= to_unsigned(integer(my_rom(511)),16);
when x"200" => lut_sig <= to_unsigned(integer(my_rom(512)),16);
when x"201" => lut_sig <= to_unsigned(integer(my_rom(513)),16);
when x"202" => lut_sig <= to_unsigned(integer(my_rom(514)),16);
when x"203" => lut_sig <= to_unsigned(integer(my_rom(515)),16);
when x"204" => lut_sig <= to_unsigned(integer(my_rom(516)),16);
when x"205" => lut_sig <= to_unsigned(integer(my_rom(517)),16);
when x"206" => lut_sig <= to_unsigned(integer(my_rom(518)),16);
when x"207" => lut_sig <= to_unsigned(integer(my_rom(519)),16);
when x"208" => lut_sig <= to_unsigned(integer(my_rom(520)),16);
when x"209" => lut_sig <= to_unsigned(integer(my_rom(521)),16);
when x"20a" => lut_sig <= to_unsigned(integer(my_rom(522)),16);
when x"20b" => lut_sig <= to_unsigned(integer(my_rom(523)),16);
when x"20c" => lut_sig <= to_unsigned(integer(my_rom(524)),16);
when x"20d" => lut_sig <= to_unsigned(integer(my_rom(525)),16);
when x"20e" => lut_sig <= to_unsigned(integer(my_rom(526)),16);
when x"20f" => lut_sig <= to_unsigned(integer(my_rom(527)),16);
when x"210" => lut_sig <= to_unsigned(integer(my_rom(528)),16);
when x"211" => lut_sig <= to_unsigned(integer(my_rom(529)),16);
when x"212" => lut_sig <= to_unsigned(integer(my_rom(530)),16);
when x"213" => lut_sig <= to_unsigned(integer(my_rom(531)),16);
when x"214" => lut_sig <= to_unsigned(integer(my_rom(532)),16);
when x"215" => lut_sig <= to_unsigned(integer(my_rom(533)),16);
when x"216" => lut_sig <= to_unsigned(integer(my_rom(534)),16);
when x"217" => lut_sig <= to_unsigned(integer(my_rom(535)),16);
when x"218" => lut_sig <= to_unsigned(integer(my_rom(536)),16);
when x"219" => lut_sig <= to_unsigned(integer(my_rom(537)),16);
when x"21a" => lut_sig <= to_unsigned(integer(my_rom(538)),16);
when x"21b" => lut_sig <= to_unsigned(integer(my_rom(539)),16);
when x"21c" => lut_sig <= to_unsigned(integer(my_rom(540)),16);
when x"21d" => lut_sig <= to_unsigned(integer(my_rom(541)),16);
when x"21e" => lut_sig <= to_unsigned(integer(my_rom(542)),16);
when x"21f" => lut_sig <= to_unsigned(integer(my_rom(543)),16);
when x"220" => lut_sig <= to_unsigned(integer(my_rom(544)),16);
when x"221" => lut_sig <= to_unsigned(integer(my_rom(545)),16);
when x"222" => lut_sig <= to_unsigned(integer(my_rom(546)),16);
when x"223" => lut_sig <= to_unsigned(integer(my_rom(547)),16);
when x"224" => lut_sig <= to_unsigned(integer(my_rom(548)),16);
when x"225" => lut_sig <= to_unsigned(integer(my_rom(549)),16);
when x"226" => lut_sig <= to_unsigned(integer(my_rom(550)),16);
when x"227" => lut_sig <= to_unsigned(integer(my_rom(551)),16);
when x"228" => lut_sig <= to_unsigned(integer(my_rom(552)),16);
when x"229" => lut_sig <= to_unsigned(integer(my_rom(553)),16);
when x"22a" => lut_sig <= to_unsigned(integer(my_rom(554)),16);
when x"22b" => lut_sig <= to_unsigned(integer(my_rom(555)),16);
when x"22c" => lut_sig <= to_unsigned(integer(my_rom(556)),16);
when x"22d" => lut_sig <= to_unsigned(integer(my_rom(557)),16);
when x"22e" => lut_sig <= to_unsigned(integer(my_rom(558)),16);
when x"22f" => lut_sig <= to_unsigned(integer(my_rom(559)),16);
when x"230" => lut_sig <= to_unsigned(integer(my_rom(560)),16);
when x"231" => lut_sig <= to_unsigned(integer(my_rom(561)),16);
when x"232" => lut_sig <= to_unsigned(integer(my_rom(562)),16);
when x"233" => lut_sig <= to_unsigned(integer(my_rom(563)),16);
when x"234" => lut_sig <= to_unsigned(integer(my_rom(564)),16);
when x"235" => lut_sig <= to_unsigned(integer(my_rom(565)),16);
when x"236" => lut_sig <= to_unsigned(integer(my_rom(566)),16);
when x"237" => lut_sig <= to_unsigned(integer(my_rom(567)),16);
when x"238" => lut_sig <= to_unsigned(integer(my_rom(568)),16);
when x"239" => lut_sig <= to_unsigned(integer(my_rom(569)),16);
when x"23a" => lut_sig <= to_unsigned(integer(my_rom(570)),16);
when x"23b" => lut_sig <= to_unsigned(integer(my_rom(571)),16);
when x"23c" => lut_sig <= to_unsigned(integer(my_rom(572)),16);
when x"23d" => lut_sig <= to_unsigned(integer(my_rom(573)),16);
when x"23e" => lut_sig <= to_unsigned(integer(my_rom(574)),16);
when x"23f" => lut_sig <= to_unsigned(integer(my_rom(575)),16);
when x"240" => lut_sig <= to_unsigned(integer(my_rom(576)),16);
when x"241" => lut_sig <= to_unsigned(integer(my_rom(577)),16);
when x"242" => lut_sig <= to_unsigned(integer(my_rom(578)),16);
when x"243" => lut_sig <= to_unsigned(integer(my_rom(579)),16);
when x"244" => lut_sig <= to_unsigned(integer(my_rom(580)),16);
when x"245" => lut_sig <= to_unsigned(integer(my_rom(581)),16);
when x"246" => lut_sig <= to_unsigned(integer(my_rom(582)),16);
when x"247" => lut_sig <= to_unsigned(integer(my_rom(583)),16);
when x"248" => lut_sig <= to_unsigned(integer(my_rom(584)),16);
when x"249" => lut_sig <= to_unsigned(integer(my_rom(585)),16);
when x"24a" => lut_sig <= to_unsigned(integer(my_rom(586)),16);
when x"24b" => lut_sig <= to_unsigned(integer(my_rom(587)),16);
when x"24c" => lut_sig <= to_unsigned(integer(my_rom(588)),16);
when x"24d" => lut_sig <= to_unsigned(integer(my_rom(589)),16);
when x"24e" => lut_sig <= to_unsigned(integer(my_rom(590)),16);
when x"24f" => lut_sig <= to_unsigned(integer(my_rom(591)),16);
when x"250" => lut_sig <= to_unsigned(integer(my_rom(592)),16);
when x"251" => lut_sig <= to_unsigned(integer(my_rom(593)),16);
when x"252" => lut_sig <= to_unsigned(integer(my_rom(594)),16);
when x"253" => lut_sig <= to_unsigned(integer(my_rom(595)),16);
when x"254" => lut_sig <= to_unsigned(integer(my_rom(596)),16);
when x"255" => lut_sig <= to_unsigned(integer(my_rom(597)),16);
when x"256" => lut_sig <= to_unsigned(integer(my_rom(598)),16);
when x"257" => lut_sig <= to_unsigned(integer(my_rom(599)),16);
when x"258" => lut_sig <= to_unsigned(integer(my_rom(600)),16);
when x"259" => lut_sig <= to_unsigned(integer(my_rom(601)),16);
when x"25a" => lut_sig <= to_unsigned(integer(my_rom(602)),16);
when x"25b" => lut_sig <= to_unsigned(integer(my_rom(603)),16);
when x"25c" => lut_sig <= to_unsigned(integer(my_rom(604)),16);
when x"25d" => lut_sig <= to_unsigned(integer(my_rom(605)),16);
when x"25e" => lut_sig <= to_unsigned(integer(my_rom(606)),16);
when x"25f" => lut_sig <= to_unsigned(integer(my_rom(607)),16);
when x"260" => lut_sig <= to_unsigned(integer(my_rom(608)),16);
when x"261" => lut_sig <= to_unsigned(integer(my_rom(609)),16);
when x"262" => lut_sig <= to_unsigned(integer(my_rom(610)),16);
when x"263" => lut_sig <= to_unsigned(integer(my_rom(611)),16);
when x"264" => lut_sig <= to_unsigned(integer(my_rom(612)),16);
when x"265" => lut_sig <= to_unsigned(integer(my_rom(613)),16);
when x"266" => lut_sig <= to_unsigned(integer(my_rom(614)),16);
when x"267" => lut_sig <= to_unsigned(integer(my_rom(615)),16);
when x"268" => lut_sig <= to_unsigned(integer(my_rom(616)),16);
when x"269" => lut_sig <= to_unsigned(integer(my_rom(617)),16);
when x"26a" => lut_sig <= to_unsigned(integer(my_rom(618)),16);
when x"26b" => lut_sig <= to_unsigned(integer(my_rom(619)),16);
when x"26c" => lut_sig <= to_unsigned(integer(my_rom(620)),16);
when x"26d" => lut_sig <= to_unsigned(integer(my_rom(621)),16);
when x"26e" => lut_sig <= to_unsigned(integer(my_rom(622)),16);
when x"26f" => lut_sig <= to_unsigned(integer(my_rom(623)),16);
when x"270" => lut_sig <= to_unsigned(integer(my_rom(624)),16);
when x"271" => lut_sig <= to_unsigned(integer(my_rom(625)),16);
when x"272" => lut_sig <= to_unsigned(integer(my_rom(626)),16);
when x"273" => lut_sig <= to_unsigned(integer(my_rom(627)),16);
when x"274" => lut_sig <= to_unsigned(integer(my_rom(628)),16);
when x"275" => lut_sig <= to_unsigned(integer(my_rom(629)),16);
when x"276" => lut_sig <= to_unsigned(integer(my_rom(630)),16);
when x"277" => lut_sig <= to_unsigned(integer(my_rom(631)),16);
when x"278" => lut_sig <= to_unsigned(integer(my_rom(632)),16);
when x"279" => lut_sig <= to_unsigned(integer(my_rom(633)),16);
when x"27a" => lut_sig <= to_unsigned(integer(my_rom(634)),16);
when x"27b" => lut_sig <= to_unsigned(integer(my_rom(635)),16);
when x"27c" => lut_sig <= to_unsigned(integer(my_rom(636)),16);
when x"27d" => lut_sig <= to_unsigned(integer(my_rom(637)),16);
when x"27e" => lut_sig <= to_unsigned(integer(my_rom(638)),16);
when x"27f" => lut_sig <= to_unsigned(integer(my_rom(639)),16);
when x"280" => lut_sig <= to_unsigned(integer(my_rom(640)),16);
when x"281" => lut_sig <= to_unsigned(integer(my_rom(641)),16);
when x"282" => lut_sig <= to_unsigned(integer(my_rom(642)),16);
when x"283" => lut_sig <= to_unsigned(integer(my_rom(643)),16);
when x"284" => lut_sig <= to_unsigned(integer(my_rom(644)),16);
when x"285" => lut_sig <= to_unsigned(integer(my_rom(645)),16);
when x"286" => lut_sig <= to_unsigned(integer(my_rom(646)),16);
when x"287" => lut_sig <= to_unsigned(integer(my_rom(647)),16);
when x"288" => lut_sig <= to_unsigned(integer(my_rom(648)),16);
when x"289" => lut_sig <= to_unsigned(integer(my_rom(649)),16);
when x"28a" => lut_sig <= to_unsigned(integer(my_rom(650)),16);
when x"28b" => lut_sig <= to_unsigned(integer(my_rom(651)),16);
when x"28c" => lut_sig <= to_unsigned(integer(my_rom(652)),16);
when x"28d" => lut_sig <= to_unsigned(integer(my_rom(653)),16);
when x"28e" => lut_sig <= to_unsigned(integer(my_rom(654)),16);
when x"28f" => lut_sig <= to_unsigned(integer(my_rom(655)),16);
when x"290" => lut_sig <= to_unsigned(integer(my_rom(656)),16);
when x"291" => lut_sig <= to_unsigned(integer(my_rom(657)),16);
when x"292" => lut_sig <= to_unsigned(integer(my_rom(658)),16);
when x"293" => lut_sig <= to_unsigned(integer(my_rom(659)),16);
when x"294" => lut_sig <= to_unsigned(integer(my_rom(660)),16);
when x"295" => lut_sig <= to_unsigned(integer(my_rom(661)),16);
when x"296" => lut_sig <= to_unsigned(integer(my_rom(662)),16);
when x"297" => lut_sig <= to_unsigned(integer(my_rom(663)),16);
when x"298" => lut_sig <= to_unsigned(integer(my_rom(664)),16);
when x"299" => lut_sig <= to_unsigned(integer(my_rom(665)),16);
when x"29a" => lut_sig <= to_unsigned(integer(my_rom(666)),16);
when x"29b" => lut_sig <= to_unsigned(integer(my_rom(667)),16);
when x"29c" => lut_sig <= to_unsigned(integer(my_rom(668)),16);
when x"29d" => lut_sig <= to_unsigned(integer(my_rom(669)),16);
when x"29e" => lut_sig <= to_unsigned(integer(my_rom(670)),16);
when x"29f" => lut_sig <= to_unsigned(integer(my_rom(671)),16);
when x"2a0" => lut_sig <= to_unsigned(integer(my_rom(672)),16);
when x"2a1" => lut_sig <= to_unsigned(integer(my_rom(673)),16);
when x"2a2" => lut_sig <= to_unsigned(integer(my_rom(674)),16);
when x"2a3" => lut_sig <= to_unsigned(integer(my_rom(675)),16);
when x"2a4" => lut_sig <= to_unsigned(integer(my_rom(676)),16);
when x"2a5" => lut_sig <= to_unsigned(integer(my_rom(677)),16);
when x"2a6" => lut_sig <= to_unsigned(integer(my_rom(678)),16);
when x"2a7" => lut_sig <= to_unsigned(integer(my_rom(679)),16);
when x"2a8" => lut_sig <= to_unsigned(integer(my_rom(680)),16);
when x"2a9" => lut_sig <= to_unsigned(integer(my_rom(681)),16);
when x"2aa" => lut_sig <= to_unsigned(integer(my_rom(682)),16);
when x"2ab" => lut_sig <= to_unsigned(integer(my_rom(683)),16);
when x"2ac" => lut_sig <= to_unsigned(integer(my_rom(684)),16);
when x"2ad" => lut_sig <= to_unsigned(integer(my_rom(685)),16);
when x"2ae" => lut_sig <= to_unsigned(integer(my_rom(686)),16);
when x"2af" => lut_sig <= to_unsigned(integer(my_rom(687)),16);
when x"2b0" => lut_sig <= to_unsigned(integer(my_rom(688)),16);
when x"2b1" => lut_sig <= to_unsigned(integer(my_rom(689)),16);
when x"2b2" => lut_sig <= to_unsigned(integer(my_rom(690)),16);
when x"2b3" => lut_sig <= to_unsigned(integer(my_rom(691)),16);
when x"2b4" => lut_sig <= to_unsigned(integer(my_rom(692)),16);
when x"2b5" => lut_sig <= to_unsigned(integer(my_rom(693)),16);
when x"2b6" => lut_sig <= to_unsigned(integer(my_rom(694)),16);
when x"2b7" => lut_sig <= to_unsigned(integer(my_rom(695)),16);
when x"2b8" => lut_sig <= to_unsigned(integer(my_rom(696)),16);
when x"2b9" => lut_sig <= to_unsigned(integer(my_rom(697)),16);
when x"2ba" => lut_sig <= to_unsigned(integer(my_rom(698)),16);
when x"2bb" => lut_sig <= to_unsigned(integer(my_rom(699)),16);
when x"2bc" => lut_sig <= to_unsigned(integer(my_rom(700)),16);
when x"2bd" => lut_sig <= to_unsigned(integer(my_rom(701)),16);
when x"2be" => lut_sig <= to_unsigned(integer(my_rom(702)),16);
when x"2bf" => lut_sig <= to_unsigned(integer(my_rom(703)),16);
when x"2c0" => lut_sig <= to_unsigned(integer(my_rom(704)),16);
when x"2c1" => lut_sig <= to_unsigned(integer(my_rom(705)),16);
when x"2c2" => lut_sig <= to_unsigned(integer(my_rom(706)),16);
when x"2c3" => lut_sig <= to_unsigned(integer(my_rom(707)),16);
when x"2c4" => lut_sig <= to_unsigned(integer(my_rom(708)),16);
when x"2c5" => lut_sig <= to_unsigned(integer(my_rom(709)),16);
when x"2c6" => lut_sig <= to_unsigned(integer(my_rom(710)),16);
when x"2c7" => lut_sig <= to_unsigned(integer(my_rom(711)),16);
when x"2c8" => lut_sig <= to_unsigned(integer(my_rom(712)),16);
when x"2c9" => lut_sig <= to_unsigned(integer(my_rom(713)),16);
when x"2ca" => lut_sig <= to_unsigned(integer(my_rom(714)),16);
when x"2cb" => lut_sig <= to_unsigned(integer(my_rom(715)),16);
when x"2cc" => lut_sig <= to_unsigned(integer(my_rom(716)),16);
when x"2cd" => lut_sig <= to_unsigned(integer(my_rom(717)),16);
when x"2ce" => lut_sig <= to_unsigned(integer(my_rom(718)),16);
when x"2cf" => lut_sig <= to_unsigned(integer(my_rom(719)),16);
when x"2d0" => lut_sig <= to_unsigned(integer(my_rom(720)),16);
when x"2d1" => lut_sig <= to_unsigned(integer(my_rom(721)),16);
when x"2d2" => lut_sig <= to_unsigned(integer(my_rom(722)),16);
when x"2d3" => lut_sig <= to_unsigned(integer(my_rom(723)),16);
when x"2d4" => lut_sig <= to_unsigned(integer(my_rom(724)),16);
when x"2d5" => lut_sig <= to_unsigned(integer(my_rom(725)),16);
when x"2d6" => lut_sig <= to_unsigned(integer(my_rom(726)),16);
when x"2d7" => lut_sig <= to_unsigned(integer(my_rom(727)),16);
when x"2d8" => lut_sig <= to_unsigned(integer(my_rom(728)),16);
when x"2d9" => lut_sig <= to_unsigned(integer(my_rom(729)),16);
when x"2da" => lut_sig <= to_unsigned(integer(my_rom(730)),16);
when x"2db" => lut_sig <= to_unsigned(integer(my_rom(731)),16);
when x"2dc" => lut_sig <= to_unsigned(integer(my_rom(732)),16);
when x"2dd" => lut_sig <= to_unsigned(integer(my_rom(733)),16);
when x"2de" => lut_sig <= to_unsigned(integer(my_rom(734)),16);
when x"2df" => lut_sig <= to_unsigned(integer(my_rom(735)),16);
when x"2e0" => lut_sig <= to_unsigned(integer(my_rom(736)),16);
when x"2e1" => lut_sig <= to_unsigned(integer(my_rom(737)),16);
when x"2e2" => lut_sig <= to_unsigned(integer(my_rom(738)),16);
when x"2e3" => lut_sig <= to_unsigned(integer(my_rom(739)),16);
when x"2e4" => lut_sig <= to_unsigned(integer(my_rom(740)),16);
when x"2e5" => lut_sig <= to_unsigned(integer(my_rom(741)),16);
when x"2e6" => lut_sig <= to_unsigned(integer(my_rom(742)),16);
when x"2e7" => lut_sig <= to_unsigned(integer(my_rom(743)),16);
when x"2e8" => lut_sig <= to_unsigned(integer(my_rom(744)),16);
when x"2e9" => lut_sig <= to_unsigned(integer(my_rom(745)),16);
when x"2ea" => lut_sig <= to_unsigned(integer(my_rom(746)),16);
when x"2eb" => lut_sig <= to_unsigned(integer(my_rom(747)),16);
when x"2ec" => lut_sig <= to_unsigned(integer(my_rom(748)),16);
when x"2ed" => lut_sig <= to_unsigned(integer(my_rom(749)),16);
when x"2ee" => lut_sig <= to_unsigned(integer(my_rom(750)),16);
when x"2ef" => lut_sig <= to_unsigned(integer(my_rom(751)),16);
when x"2f0" => lut_sig <= to_unsigned(integer(my_rom(752)),16);
when x"2f1" => lut_sig <= to_unsigned(integer(my_rom(753)),16);
when x"2f2" => lut_sig <= to_unsigned(integer(my_rom(754)),16);
when x"2f3" => lut_sig <= to_unsigned(integer(my_rom(755)),16);
when x"2f4" => lut_sig <= to_unsigned(integer(my_rom(756)),16);
when x"2f5" => lut_sig <= to_unsigned(integer(my_rom(757)),16);
when x"2f6" => lut_sig <= to_unsigned(integer(my_rom(758)),16);
when x"2f7" => lut_sig <= to_unsigned(integer(my_rom(759)),16);
when x"2f8" => lut_sig <= to_unsigned(integer(my_rom(760)),16);
when x"2f9" => lut_sig <= to_unsigned(integer(my_rom(761)),16);
when x"2fa" => lut_sig <= to_unsigned(integer(my_rom(762)),16);
when x"2fb" => lut_sig <= to_unsigned(integer(my_rom(763)),16);
when x"2fc" => lut_sig <= to_unsigned(integer(my_rom(764)),16);
when x"2fd" => lut_sig <= to_unsigned(integer(my_rom(765)),16);
when x"2fe" => lut_sig <= to_unsigned(integer(my_rom(766)),16);
when x"2ff" => lut_sig <= to_unsigned(integer(my_rom(767)),16);
when x"300" => lut_sig <= to_unsigned(integer(my_rom(768)),16);
when x"301" => lut_sig <= to_unsigned(integer(my_rom(769)),16);
when x"302" => lut_sig <= to_unsigned(integer(my_rom(770)),16);
when x"303" => lut_sig <= to_unsigned(integer(my_rom(771)),16);
when x"304" => lut_sig <= to_unsigned(integer(my_rom(772)),16);
when x"305" => lut_sig <= to_unsigned(integer(my_rom(773)),16);
when x"306" => lut_sig <= to_unsigned(integer(my_rom(774)),16);
when x"307" => lut_sig <= to_unsigned(integer(my_rom(775)),16);
when x"308" => lut_sig <= to_unsigned(integer(my_rom(776)),16);
when x"309" => lut_sig <= to_unsigned(integer(my_rom(777)),16);
when x"30a" => lut_sig <= to_unsigned(integer(my_rom(778)),16);
when x"30b" => lut_sig <= to_unsigned(integer(my_rom(779)),16);
when x"30c" => lut_sig <= to_unsigned(integer(my_rom(780)),16);
when x"30d" => lut_sig <= to_unsigned(integer(my_rom(781)),16);
when x"30e" => lut_sig <= to_unsigned(integer(my_rom(782)),16);
when x"30f" => lut_sig <= to_unsigned(integer(my_rom(783)),16);
when x"310" => lut_sig <= to_unsigned(integer(my_rom(784)),16);
when x"311" => lut_sig <= to_unsigned(integer(my_rom(785)),16);
when x"312" => lut_sig <= to_unsigned(integer(my_rom(786)),16);
when x"313" => lut_sig <= to_unsigned(integer(my_rom(787)),16);
when x"314" => lut_sig <= to_unsigned(integer(my_rom(788)),16);
when x"315" => lut_sig <= to_unsigned(integer(my_rom(789)),16);
when x"316" => lut_sig <= to_unsigned(integer(my_rom(790)),16);
when x"317" => lut_sig <= to_unsigned(integer(my_rom(791)),16);
when x"318" => lut_sig <= to_unsigned(integer(my_rom(792)),16);
when x"319" => lut_sig <= to_unsigned(integer(my_rom(793)),16);
when x"31a" => lut_sig <= to_unsigned(integer(my_rom(794)),16);
when x"31b" => lut_sig <= to_unsigned(integer(my_rom(795)),16);
when x"31c" => lut_sig <= to_unsigned(integer(my_rom(796)),16);
when x"31d" => lut_sig <= to_unsigned(integer(my_rom(797)),16);
when x"31e" => lut_sig <= to_unsigned(integer(my_rom(798)),16);
when x"31f" => lut_sig <= to_unsigned(integer(my_rom(799)),16);
when x"320" => lut_sig <= to_unsigned(integer(my_rom(800)),16);
when x"321" => lut_sig <= to_unsigned(integer(my_rom(801)),16);
when x"322" => lut_sig <= to_unsigned(integer(my_rom(802)),16);
when x"323" => lut_sig <= to_unsigned(integer(my_rom(803)),16);
when x"324" => lut_sig <= to_unsigned(integer(my_rom(804)),16);
when x"325" => lut_sig <= to_unsigned(integer(my_rom(805)),16);
when x"326" => lut_sig <= to_unsigned(integer(my_rom(806)),16);
when x"327" => lut_sig <= to_unsigned(integer(my_rom(807)),16);
when x"328" => lut_sig <= to_unsigned(integer(my_rom(808)),16);
when x"329" => lut_sig <= to_unsigned(integer(my_rom(809)),16);
when x"32a" => lut_sig <= to_unsigned(integer(my_rom(810)),16);
when x"32b" => lut_sig <= to_unsigned(integer(my_rom(811)),16);
when x"32c" => lut_sig <= to_unsigned(integer(my_rom(812)),16);
when x"32d" => lut_sig <= to_unsigned(integer(my_rom(813)),16);
when x"32e" => lut_sig <= to_unsigned(integer(my_rom(814)),16);
when x"32f" => lut_sig <= to_unsigned(integer(my_rom(815)),16);
when x"330" => lut_sig <= to_unsigned(integer(my_rom(816)),16);
when x"331" => lut_sig <= to_unsigned(integer(my_rom(817)),16);
when x"332" => lut_sig <= to_unsigned(integer(my_rom(818)),16);
when x"333" => lut_sig <= to_unsigned(integer(my_rom(819)),16);
when x"334" => lut_sig <= to_unsigned(integer(my_rom(820)),16);
when x"335" => lut_sig <= to_unsigned(integer(my_rom(821)),16);
when x"336" => lut_sig <= to_unsigned(integer(my_rom(822)),16);
when x"337" => lut_sig <= to_unsigned(integer(my_rom(823)),16);
when x"338" => lut_sig <= to_unsigned(integer(my_rom(824)),16);
when x"339" => lut_sig <= to_unsigned(integer(my_rom(825)),16);
when x"33a" => lut_sig <= to_unsigned(integer(my_rom(826)),16);
when x"33b" => lut_sig <= to_unsigned(integer(my_rom(827)),16);
when x"33c" => lut_sig <= to_unsigned(integer(my_rom(828)),16);
when x"33d" => lut_sig <= to_unsigned(integer(my_rom(829)),16);
when x"33e" => lut_sig <= to_unsigned(integer(my_rom(830)),16);
when x"33f" => lut_sig <= to_unsigned(integer(my_rom(831)),16);
when x"340" => lut_sig <= to_unsigned(integer(my_rom(832)),16);
when x"341" => lut_sig <= to_unsigned(integer(my_rom(833)),16);
when x"342" => lut_sig <= to_unsigned(integer(my_rom(834)),16);
when x"343" => lut_sig <= to_unsigned(integer(my_rom(835)),16);
when x"344" => lut_sig <= to_unsigned(integer(my_rom(836)),16);
when x"345" => lut_sig <= to_unsigned(integer(my_rom(837)),16);
when x"346" => lut_sig <= to_unsigned(integer(my_rom(838)),16);
when x"347" => lut_sig <= to_unsigned(integer(my_rom(839)),16);
when x"348" => lut_sig <= to_unsigned(integer(my_rom(840)),16);
when x"349" => lut_sig <= to_unsigned(integer(my_rom(841)),16);
when x"34a" => lut_sig <= to_unsigned(integer(my_rom(842)),16);
when x"34b" => lut_sig <= to_unsigned(integer(my_rom(843)),16);
when x"34c" => lut_sig <= to_unsigned(integer(my_rom(844)),16);
when x"34d" => lut_sig <= to_unsigned(integer(my_rom(845)),16);
when x"34e" => lut_sig <= to_unsigned(integer(my_rom(846)),16);
when x"34f" => lut_sig <= to_unsigned(integer(my_rom(847)),16);
when x"350" => lut_sig <= to_unsigned(integer(my_rom(848)),16);
when x"351" => lut_sig <= to_unsigned(integer(my_rom(849)),16);
when x"352" => lut_sig <= to_unsigned(integer(my_rom(850)),16);
when x"353" => lut_sig <= to_unsigned(integer(my_rom(851)),16);
when x"354" => lut_sig <= to_unsigned(integer(my_rom(852)),16);
when x"355" => lut_sig <= to_unsigned(integer(my_rom(853)),16);
when x"356" => lut_sig <= to_unsigned(integer(my_rom(854)),16);
when x"357" => lut_sig <= to_unsigned(integer(my_rom(855)),16);
when x"358" => lut_sig <= to_unsigned(integer(my_rom(856)),16);
when x"359" => lut_sig <= to_unsigned(integer(my_rom(857)),16);
when x"35a" => lut_sig <= to_unsigned(integer(my_rom(858)),16);
when x"35b" => lut_sig <= to_unsigned(integer(my_rom(859)),16);
when x"35c" => lut_sig <= to_unsigned(integer(my_rom(860)),16);
when x"35d" => lut_sig <= to_unsigned(integer(my_rom(861)),16);
when x"35e" => lut_sig <= to_unsigned(integer(my_rom(862)),16);
when x"35f" => lut_sig <= to_unsigned(integer(my_rom(863)),16);
when x"360" => lut_sig <= to_unsigned(integer(my_rom(864)),16);
when x"361" => lut_sig <= to_unsigned(integer(my_rom(865)),16);
when x"362" => lut_sig <= to_unsigned(integer(my_rom(866)),16);
when x"363" => lut_sig <= to_unsigned(integer(my_rom(867)),16);
when x"364" => lut_sig <= to_unsigned(integer(my_rom(868)),16);
when x"365" => lut_sig <= to_unsigned(integer(my_rom(869)),16);
when x"366" => lut_sig <= to_unsigned(integer(my_rom(870)),16);
when x"367" => lut_sig <= to_unsigned(integer(my_rom(871)),16);
when x"368" => lut_sig <= to_unsigned(integer(my_rom(872)),16);
when x"369" => lut_sig <= to_unsigned(integer(my_rom(873)),16);
when x"36a" => lut_sig <= to_unsigned(integer(my_rom(874)),16);
when x"36b" => lut_sig <= to_unsigned(integer(my_rom(875)),16);
when x"36c" => lut_sig <= to_unsigned(integer(my_rom(876)),16);
when x"36d" => lut_sig <= to_unsigned(integer(my_rom(877)),16);
when x"36e" => lut_sig <= to_unsigned(integer(my_rom(878)),16);
when x"36f" => lut_sig <= to_unsigned(integer(my_rom(879)),16);
when x"370" => lut_sig <= to_unsigned(integer(my_rom(880)),16);
when x"371" => lut_sig <= to_unsigned(integer(my_rom(881)),16);
when x"372" => lut_sig <= to_unsigned(integer(my_rom(882)),16);
when x"373" => lut_sig <= to_unsigned(integer(my_rom(883)),16);
when x"374" => lut_sig <= to_unsigned(integer(my_rom(884)),16);
when x"375" => lut_sig <= to_unsigned(integer(my_rom(885)),16);
when x"376" => lut_sig <= to_unsigned(integer(my_rom(886)),16);
when x"377" => lut_sig <= to_unsigned(integer(my_rom(887)),16);
when x"378" => lut_sig <= to_unsigned(integer(my_rom(888)),16);
when x"379" => lut_sig <= to_unsigned(integer(my_rom(889)),16);
when x"37a" => lut_sig <= to_unsigned(integer(my_rom(890)),16);
when x"37b" => lut_sig <= to_unsigned(integer(my_rom(891)),16);
when x"37c" => lut_sig <= to_unsigned(integer(my_rom(892)),16);
when x"37d" => lut_sig <= to_unsigned(integer(my_rom(893)),16);
when x"37e" => lut_sig <= to_unsigned(integer(my_rom(894)),16);
when x"37f" => lut_sig <= to_unsigned(integer(my_rom(895)),16);
when x"380" => lut_sig <= to_unsigned(integer(my_rom(896)),16);
when x"381" => lut_sig <= to_unsigned(integer(my_rom(897)),16);
when x"382" => lut_sig <= to_unsigned(integer(my_rom(898)),16);
when x"383" => lut_sig <= to_unsigned(integer(my_rom(899)),16);
when x"384" => lut_sig <= to_unsigned(integer(my_rom(900)),16);
when x"385" => lut_sig <= to_unsigned(integer(my_rom(901)),16);
when x"386" => lut_sig <= to_unsigned(integer(my_rom(902)),16);
when x"387" => lut_sig <= to_unsigned(integer(my_rom(903)),16);
when x"388" => lut_sig <= to_unsigned(integer(my_rom(904)),16);
when x"389" => lut_sig <= to_unsigned(integer(my_rom(905)),16);
when x"38a" => lut_sig <= to_unsigned(integer(my_rom(906)),16);
when x"38b" => lut_sig <= to_unsigned(integer(my_rom(907)),16);
when x"38c" => lut_sig <= to_unsigned(integer(my_rom(908)),16);
when x"38d" => lut_sig <= to_unsigned(integer(my_rom(909)),16);
when x"38e" => lut_sig <= to_unsigned(integer(my_rom(910)),16);
when x"38f" => lut_sig <= to_unsigned(integer(my_rom(911)),16);
when x"390" => lut_sig <= to_unsigned(integer(my_rom(912)),16);
when x"391" => lut_sig <= to_unsigned(integer(my_rom(913)),16);
when x"392" => lut_sig <= to_unsigned(integer(my_rom(914)),16);
when x"393" => lut_sig <= to_unsigned(integer(my_rom(915)),16);
when x"394" => lut_sig <= to_unsigned(integer(my_rom(916)),16);
when x"395" => lut_sig <= to_unsigned(integer(my_rom(917)),16);
when x"396" => lut_sig <= to_unsigned(integer(my_rom(918)),16);
when x"397" => lut_sig <= to_unsigned(integer(my_rom(919)),16);
when x"398" => lut_sig <= to_unsigned(integer(my_rom(920)),16);
when x"399" => lut_sig <= to_unsigned(integer(my_rom(921)),16);
when x"39a" => lut_sig <= to_unsigned(integer(my_rom(922)),16);
when x"39b" => lut_sig <= to_unsigned(integer(my_rom(923)),16);
when x"39c" => lut_sig <= to_unsigned(integer(my_rom(924)),16);
when x"39d" => lut_sig <= to_unsigned(integer(my_rom(925)),16);
when x"39e" => lut_sig <= to_unsigned(integer(my_rom(926)),16);
when x"39f" => lut_sig <= to_unsigned(integer(my_rom(927)),16);
when x"3a0" => lut_sig <= to_unsigned(integer(my_rom(928)),16);
when x"3a1" => lut_sig <= to_unsigned(integer(my_rom(929)),16);
when x"3a2" => lut_sig <= to_unsigned(integer(my_rom(930)),16);
when x"3a3" => lut_sig <= to_unsigned(integer(my_rom(931)),16);
when x"3a4" => lut_sig <= to_unsigned(integer(my_rom(932)),16);
when x"3a5" => lut_sig <= to_unsigned(integer(my_rom(933)),16);
when x"3a6" => lut_sig <= to_unsigned(integer(my_rom(934)),16);
when x"3a7" => lut_sig <= to_unsigned(integer(my_rom(935)),16);
when x"3a8" => lut_sig <= to_unsigned(integer(my_rom(936)),16);
when x"3a9" => lut_sig <= to_unsigned(integer(my_rom(937)),16);
when x"3aa" => lut_sig <= to_unsigned(integer(my_rom(938)),16);
when x"3ab" => lut_sig <= to_unsigned(integer(my_rom(939)),16);
when x"3ac" => lut_sig <= to_unsigned(integer(my_rom(940)),16);
when x"3ad" => lut_sig <= to_unsigned(integer(my_rom(941)),16);
when x"3ae" => lut_sig <= to_unsigned(integer(my_rom(942)),16);
when x"3af" => lut_sig <= to_unsigned(integer(my_rom(943)),16);
when x"3b0" => lut_sig <= to_unsigned(integer(my_rom(944)),16);
when x"3b1" => lut_sig <= to_unsigned(integer(my_rom(945)),16);
when x"3b2" => lut_sig <= to_unsigned(integer(my_rom(946)),16);
when x"3b3" => lut_sig <= to_unsigned(integer(my_rom(947)),16);
when x"3b4" => lut_sig <= to_unsigned(integer(my_rom(948)),16);
when x"3b5" => lut_sig <= to_unsigned(integer(my_rom(949)),16);
when x"3b6" => lut_sig <= to_unsigned(integer(my_rom(950)),16);
when x"3b7" => lut_sig <= to_unsigned(integer(my_rom(951)),16);
when x"3b8" => lut_sig <= to_unsigned(integer(my_rom(952)),16);
when x"3b9" => lut_sig <= to_unsigned(integer(my_rom(953)),16);
when x"3ba" => lut_sig <= to_unsigned(integer(my_rom(954)),16);
when x"3bb" => lut_sig <= to_unsigned(integer(my_rom(955)),16);
when x"3bc" => lut_sig <= to_unsigned(integer(my_rom(956)),16);
when x"3bd" => lut_sig <= to_unsigned(integer(my_rom(957)),16);
when x"3be" => lut_sig <= to_unsigned(integer(my_rom(958)),16);
when x"3bf" => lut_sig <= to_unsigned(integer(my_rom(959)),16);
when x"3c0" => lut_sig <= to_unsigned(integer(my_rom(960)),16);
when x"3c1" => lut_sig <= to_unsigned(integer(my_rom(961)),16);
when x"3c2" => lut_sig <= to_unsigned(integer(my_rom(962)),16);
when x"3c3" => lut_sig <= to_unsigned(integer(my_rom(963)),16);
when x"3c4" => lut_sig <= to_unsigned(integer(my_rom(964)),16);
when x"3c5" => lut_sig <= to_unsigned(integer(my_rom(965)),16);
when x"3c6" => lut_sig <= to_unsigned(integer(my_rom(966)),16);
when x"3c7" => lut_sig <= to_unsigned(integer(my_rom(967)),16);
when x"3c8" => lut_sig <= to_unsigned(integer(my_rom(968)),16);
when x"3c9" => lut_sig <= to_unsigned(integer(my_rom(969)),16);
when x"3ca" => lut_sig <= to_unsigned(integer(my_rom(970)),16);
when x"3cb" => lut_sig <= to_unsigned(integer(my_rom(971)),16);
when x"3cc" => lut_sig <= to_unsigned(integer(my_rom(972)),16);
when x"3cd" => lut_sig <= to_unsigned(integer(my_rom(973)),16);
when x"3ce" => lut_sig <= to_unsigned(integer(my_rom(974)),16);
when x"3cf" => lut_sig <= to_unsigned(integer(my_rom(975)),16);
when x"3d0" => lut_sig <= to_unsigned(integer(my_rom(976)),16);
when x"3d1" => lut_sig <= to_unsigned(integer(my_rom(977)),16);
when x"3d2" => lut_sig <= to_unsigned(integer(my_rom(978)),16);
when x"3d3" => lut_sig <= to_unsigned(integer(my_rom(979)),16);
when x"3d4" => lut_sig <= to_unsigned(integer(my_rom(980)),16);
when x"3d5" => lut_sig <= to_unsigned(integer(my_rom(981)),16);
when x"3d6" => lut_sig <= to_unsigned(integer(my_rom(982)),16);
when x"3d7" => lut_sig <= to_unsigned(integer(my_rom(983)),16);
when x"3d8" => lut_sig <= to_unsigned(integer(my_rom(984)),16);
when x"3d9" => lut_sig <= to_unsigned(integer(my_rom(985)),16);
when x"3da" => lut_sig <= to_unsigned(integer(my_rom(986)),16);
when x"3db" => lut_sig <= to_unsigned(integer(my_rom(987)),16);
when x"3dc" => lut_sig <= to_unsigned(integer(my_rom(988)),16);
when x"3dd" => lut_sig <= to_unsigned(integer(my_rom(989)),16);
when x"3de" => lut_sig <= to_unsigned(integer(my_rom(990)),16);
when x"3df" => lut_sig <= to_unsigned(integer(my_rom(991)),16);
when x"3e0" => lut_sig <= to_unsigned(integer(my_rom(992)),16);
when x"3e1" => lut_sig <= to_unsigned(integer(my_rom(993)),16);
when x"3e2" => lut_sig <= to_unsigned(integer(my_rom(994)),16);
when x"3e3" => lut_sig <= to_unsigned(integer(my_rom(995)),16);
when x"3e4" => lut_sig <= to_unsigned(integer(my_rom(996)),16);
when x"3e5" => lut_sig <= to_unsigned(integer(my_rom(997)),16);
when x"3e6" => lut_sig <= to_unsigned(integer(my_rom(998)),16);
when x"3e7" => lut_sig <= to_unsigned(integer(my_rom(999)),16);
when x"3e8" => lut_sig <= to_unsigned(integer(my_rom(1000)),16);
when x"3e9" => lut_sig <= to_unsigned(integer(my_rom(1001)),16);
when x"3ea" => lut_sig <= to_unsigned(integer(my_rom(1002)),16);
when x"3eb" => lut_sig <= to_unsigned(integer(my_rom(1003)),16);
when x"3ec" => lut_sig <= to_unsigned(integer(my_rom(1004)),16);
when x"3ed" => lut_sig <= to_unsigned(integer(my_rom(1005)),16);
when x"3ee" => lut_sig <= to_unsigned(integer(my_rom(1006)),16);
when x"3ef" => lut_sig <= to_unsigned(integer(my_rom(1007)),16);
when x"3f0" => lut_sig <= to_unsigned(integer(my_rom(1008)),16);
when x"3f1" => lut_sig <= to_unsigned(integer(my_rom(1009)),16);
when x"3f2" => lut_sig <= to_unsigned(integer(my_rom(1010)),16);
when x"3f3" => lut_sig <= to_unsigned(integer(my_rom(1011)),16);
when x"3f4" => lut_sig <= to_unsigned(integer(my_rom(1012)),16);
when x"3f5" => lut_sig <= to_unsigned(integer(my_rom(1013)),16);
when x"3f6" => lut_sig <= to_unsigned(integer(my_rom(1014)),16);
when x"3f7" => lut_sig <= to_unsigned(integer(my_rom(1015)),16);
when x"3f8" => lut_sig <= to_unsigned(integer(my_rom(1016)),16);
when x"3f9" => lut_sig <= to_unsigned(integer(my_rom(1017)),16);
when x"3fa" => lut_sig <= to_unsigned(integer(my_rom(1018)),16);
when x"3fb" => lut_sig <= to_unsigned(integer(my_rom(1019)),16);
when x"3fc" => lut_sig <= to_unsigned(integer(my_rom(1020)),16);
when x"3fd" => lut_sig <= to_unsigned(integer(my_rom(1021)),16);
when x"3fe" => lut_sig <= to_unsigned(integer(my_rom(1022)),16);
when x"3ff" => lut_sig <= to_unsigned(integer(my_rom(1023)),16);
when x"400" => lut_sig <= to_unsigned(integer(my_rom(1024)),16);
when x"401" => lut_sig <= to_unsigned(integer(my_rom(1025)),16);
when x"402" => lut_sig <= to_unsigned(integer(my_rom(1026)),16);
when x"403" => lut_sig <= to_unsigned(integer(my_rom(1027)),16);
when x"404" => lut_sig <= to_unsigned(integer(my_rom(1028)),16);
when x"405" => lut_sig <= to_unsigned(integer(my_rom(1029)),16);
when x"406" => lut_sig <= to_unsigned(integer(my_rom(1030)),16);
when x"407" => lut_sig <= to_unsigned(integer(my_rom(1031)),16);
when x"408" => lut_sig <= to_unsigned(integer(my_rom(1032)),16);
when x"409" => lut_sig <= to_unsigned(integer(my_rom(1033)),16);
when x"40a" => lut_sig <= to_unsigned(integer(my_rom(1034)),16);
when x"40b" => lut_sig <= to_unsigned(integer(my_rom(1035)),16);
when x"40c" => lut_sig <= to_unsigned(integer(my_rom(1036)),16);
when x"40d" => lut_sig <= to_unsigned(integer(my_rom(1037)),16);
when x"40e" => lut_sig <= to_unsigned(integer(my_rom(1038)),16);
when x"40f" => lut_sig <= to_unsigned(integer(my_rom(1039)),16);
when x"410" => lut_sig <= to_unsigned(integer(my_rom(1040)),16);
when x"411" => lut_sig <= to_unsigned(integer(my_rom(1041)),16);
when x"412" => lut_sig <= to_unsigned(integer(my_rom(1042)),16);
when x"413" => lut_sig <= to_unsigned(integer(my_rom(1043)),16);
when x"414" => lut_sig <= to_unsigned(integer(my_rom(1044)),16);
when x"415" => lut_sig <= to_unsigned(integer(my_rom(1045)),16);
when x"416" => lut_sig <= to_unsigned(integer(my_rom(1046)),16);
when x"417" => lut_sig <= to_unsigned(integer(my_rom(1047)),16);
when x"418" => lut_sig <= to_unsigned(integer(my_rom(1048)),16);
when x"419" => lut_sig <= to_unsigned(integer(my_rom(1049)),16);
when x"41a" => lut_sig <= to_unsigned(integer(my_rom(1050)),16);
when x"41b" => lut_sig <= to_unsigned(integer(my_rom(1051)),16);
when x"41c" => lut_sig <= to_unsigned(integer(my_rom(1052)),16);
when x"41d" => lut_sig <= to_unsigned(integer(my_rom(1053)),16);
when x"41e" => lut_sig <= to_unsigned(integer(my_rom(1054)),16);
when x"41f" => lut_sig <= to_unsigned(integer(my_rom(1055)),16);
when x"420" => lut_sig <= to_unsigned(integer(my_rom(1056)),16);
when x"421" => lut_sig <= to_unsigned(integer(my_rom(1057)),16);
when x"422" => lut_sig <= to_unsigned(integer(my_rom(1058)),16);
when x"423" => lut_sig <= to_unsigned(integer(my_rom(1059)),16);
when x"424" => lut_sig <= to_unsigned(integer(my_rom(1060)),16);
when x"425" => lut_sig <= to_unsigned(integer(my_rom(1061)),16);
when x"426" => lut_sig <= to_unsigned(integer(my_rom(1062)),16);
when x"427" => lut_sig <= to_unsigned(integer(my_rom(1063)),16);
when x"428" => lut_sig <= to_unsigned(integer(my_rom(1064)),16);
when x"429" => lut_sig <= to_unsigned(integer(my_rom(1065)),16);
when x"42a" => lut_sig <= to_unsigned(integer(my_rom(1066)),16);
when x"42b" => lut_sig <= to_unsigned(integer(my_rom(1067)),16);
when x"42c" => lut_sig <= to_unsigned(integer(my_rom(1068)),16);
when x"42d" => lut_sig <= to_unsigned(integer(my_rom(1069)),16);
when x"42e" => lut_sig <= to_unsigned(integer(my_rom(1070)),16);
when x"42f" => lut_sig <= to_unsigned(integer(my_rom(1071)),16);
when x"430" => lut_sig <= to_unsigned(integer(my_rom(1072)),16);
when x"431" => lut_sig <= to_unsigned(integer(my_rom(1073)),16);
when x"432" => lut_sig <= to_unsigned(integer(my_rom(1074)),16);
when x"433" => lut_sig <= to_unsigned(integer(my_rom(1075)),16);
when x"434" => lut_sig <= to_unsigned(integer(my_rom(1076)),16);
when x"435" => lut_sig <= to_unsigned(integer(my_rom(1077)),16);
when x"436" => lut_sig <= to_unsigned(integer(my_rom(1078)),16);
when x"437" => lut_sig <= to_unsigned(integer(my_rom(1079)),16);
when x"438" => lut_sig <= to_unsigned(integer(my_rom(1080)),16);
when x"439" => lut_sig <= to_unsigned(integer(my_rom(1081)),16);
when x"43a" => lut_sig <= to_unsigned(integer(my_rom(1082)),16);
when x"43b" => lut_sig <= to_unsigned(integer(my_rom(1083)),16);
when x"43c" => lut_sig <= to_unsigned(integer(my_rom(1084)),16);
when x"43d" => lut_sig <= to_unsigned(integer(my_rom(1085)),16);
when x"43e" => lut_sig <= to_unsigned(integer(my_rom(1086)),16);
when x"43f" => lut_sig <= to_unsigned(integer(my_rom(1087)),16);
when x"440" => lut_sig <= to_unsigned(integer(my_rom(1088)),16);
when x"441" => lut_sig <= to_unsigned(integer(my_rom(1089)),16);
when x"442" => lut_sig <= to_unsigned(integer(my_rom(1090)),16);
when x"443" => lut_sig <= to_unsigned(integer(my_rom(1091)),16);
when x"444" => lut_sig <= to_unsigned(integer(my_rom(1092)),16);
when x"445" => lut_sig <= to_unsigned(integer(my_rom(1093)),16);
when x"446" => lut_sig <= to_unsigned(integer(my_rom(1094)),16);
when x"447" => lut_sig <= to_unsigned(integer(my_rom(1095)),16);
when x"448" => lut_sig <= to_unsigned(integer(my_rom(1096)),16);
when x"449" => lut_sig <= to_unsigned(integer(my_rom(1097)),16);
when x"44a" => lut_sig <= to_unsigned(integer(my_rom(1098)),16);
when x"44b" => lut_sig <= to_unsigned(integer(my_rom(1099)),16);
when x"44c" => lut_sig <= to_unsigned(integer(my_rom(1100)),16);
when x"44d" => lut_sig <= to_unsigned(integer(my_rom(1101)),16);
when x"44e" => lut_sig <= to_unsigned(integer(my_rom(1102)),16);
when x"44f" => lut_sig <= to_unsigned(integer(my_rom(1103)),16);
when x"450" => lut_sig <= to_unsigned(integer(my_rom(1104)),16);
when x"451" => lut_sig <= to_unsigned(integer(my_rom(1105)),16);
when x"452" => lut_sig <= to_unsigned(integer(my_rom(1106)),16);
when x"453" => lut_sig <= to_unsigned(integer(my_rom(1107)),16);
when x"454" => lut_sig <= to_unsigned(integer(my_rom(1108)),16);
when x"455" => lut_sig <= to_unsigned(integer(my_rom(1109)),16);
when x"456" => lut_sig <= to_unsigned(integer(my_rom(1110)),16);
when x"457" => lut_sig <= to_unsigned(integer(my_rom(1111)),16);
when x"458" => lut_sig <= to_unsigned(integer(my_rom(1112)),16);
when x"459" => lut_sig <= to_unsigned(integer(my_rom(1113)),16);
when x"45a" => lut_sig <= to_unsigned(integer(my_rom(1114)),16);
when x"45b" => lut_sig <= to_unsigned(integer(my_rom(1115)),16);
when x"45c" => lut_sig <= to_unsigned(integer(my_rom(1116)),16);
when x"45d" => lut_sig <= to_unsigned(integer(my_rom(1117)),16);
when x"45e" => lut_sig <= to_unsigned(integer(my_rom(1118)),16);
when x"45f" => lut_sig <= to_unsigned(integer(my_rom(1119)),16);
when x"460" => lut_sig <= to_unsigned(integer(my_rom(1120)),16);
when x"461" => lut_sig <= to_unsigned(integer(my_rom(1121)),16);
when x"462" => lut_sig <= to_unsigned(integer(my_rom(1122)),16);
when x"463" => lut_sig <= to_unsigned(integer(my_rom(1123)),16);
when x"464" => lut_sig <= to_unsigned(integer(my_rom(1124)),16);
when x"465" => lut_sig <= to_unsigned(integer(my_rom(1125)),16);
when x"466" => lut_sig <= to_unsigned(integer(my_rom(1126)),16);
when x"467" => lut_sig <= to_unsigned(integer(my_rom(1127)),16);
when x"468" => lut_sig <= to_unsigned(integer(my_rom(1128)),16);
when x"469" => lut_sig <= to_unsigned(integer(my_rom(1129)),16);
when x"46a" => lut_sig <= to_unsigned(integer(my_rom(1130)),16);
when x"46b" => lut_sig <= to_unsigned(integer(my_rom(1131)),16);
when x"46c" => lut_sig <= to_unsigned(integer(my_rom(1132)),16);
when x"46d" => lut_sig <= to_unsigned(integer(my_rom(1133)),16);
when x"46e" => lut_sig <= to_unsigned(integer(my_rom(1134)),16);
when x"46f" => lut_sig <= to_unsigned(integer(my_rom(1135)),16);
when x"470" => lut_sig <= to_unsigned(integer(my_rom(1136)),16);
when x"471" => lut_sig <= to_unsigned(integer(my_rom(1137)),16);
when x"472" => lut_sig <= to_unsigned(integer(my_rom(1138)),16);
when x"473" => lut_sig <= to_unsigned(integer(my_rom(1139)),16);
when x"474" => lut_sig <= to_unsigned(integer(my_rom(1140)),16);
when x"475" => lut_sig <= to_unsigned(integer(my_rom(1141)),16);
when x"476" => lut_sig <= to_unsigned(integer(my_rom(1142)),16);
when x"477" => lut_sig <= to_unsigned(integer(my_rom(1143)),16);
when x"478" => lut_sig <= to_unsigned(integer(my_rom(1144)),16);
when x"479" => lut_sig <= to_unsigned(integer(my_rom(1145)),16);
when x"47a" => lut_sig <= to_unsigned(integer(my_rom(1146)),16);
when x"47b" => lut_sig <= to_unsigned(integer(my_rom(1147)),16);
when x"47c" => lut_sig <= to_unsigned(integer(my_rom(1148)),16);
when x"47d" => lut_sig <= to_unsigned(integer(my_rom(1149)),16);
when x"47e" => lut_sig <= to_unsigned(integer(my_rom(1150)),16);
when x"47f" => lut_sig <= to_unsigned(integer(my_rom(1151)),16);
when x"480" => lut_sig <= to_unsigned(integer(my_rom(1152)),16);
when x"481" => lut_sig <= to_unsigned(integer(my_rom(1153)),16);
when x"482" => lut_sig <= to_unsigned(integer(my_rom(1154)),16);
when x"483" => lut_sig <= to_unsigned(integer(my_rom(1155)),16);
when x"484" => lut_sig <= to_unsigned(integer(my_rom(1156)),16);
when x"485" => lut_sig <= to_unsigned(integer(my_rom(1157)),16);
when x"486" => lut_sig <= to_unsigned(integer(my_rom(1158)),16);
when x"487" => lut_sig <= to_unsigned(integer(my_rom(1159)),16);
when x"488" => lut_sig <= to_unsigned(integer(my_rom(1160)),16);
when x"489" => lut_sig <= to_unsigned(integer(my_rom(1161)),16);
when x"48a" => lut_sig <= to_unsigned(integer(my_rom(1162)),16);
when x"48b" => lut_sig <= to_unsigned(integer(my_rom(1163)),16);
when x"48c" => lut_sig <= to_unsigned(integer(my_rom(1164)),16);
when x"48d" => lut_sig <= to_unsigned(integer(my_rom(1165)),16);
when x"48e" => lut_sig <= to_unsigned(integer(my_rom(1166)),16);
when x"48f" => lut_sig <= to_unsigned(integer(my_rom(1167)),16);
when x"490" => lut_sig <= to_unsigned(integer(my_rom(1168)),16);
when x"491" => lut_sig <= to_unsigned(integer(my_rom(1169)),16);
when x"492" => lut_sig <= to_unsigned(integer(my_rom(1170)),16);
when x"493" => lut_sig <= to_unsigned(integer(my_rom(1171)),16);
when x"494" => lut_sig <= to_unsigned(integer(my_rom(1172)),16);
when x"495" => lut_sig <= to_unsigned(integer(my_rom(1173)),16);
when x"496" => lut_sig <= to_unsigned(integer(my_rom(1174)),16);
when x"497" => lut_sig <= to_unsigned(integer(my_rom(1175)),16);
when x"498" => lut_sig <= to_unsigned(integer(my_rom(1176)),16);
when x"499" => lut_sig <= to_unsigned(integer(my_rom(1177)),16);
when x"49a" => lut_sig <= to_unsigned(integer(my_rom(1178)),16);
when x"49b" => lut_sig <= to_unsigned(integer(my_rom(1179)),16);
when x"49c" => lut_sig <= to_unsigned(integer(my_rom(1180)),16);
when x"49d" => lut_sig <= to_unsigned(integer(my_rom(1181)),16);
when x"49e" => lut_sig <= to_unsigned(integer(my_rom(1182)),16);
when x"49f" => lut_sig <= to_unsigned(integer(my_rom(1183)),16);
when x"4a0" => lut_sig <= to_unsigned(integer(my_rom(1184)),16);
when x"4a1" => lut_sig <= to_unsigned(integer(my_rom(1185)),16);
when x"4a2" => lut_sig <= to_unsigned(integer(my_rom(1186)),16);
when x"4a3" => lut_sig <= to_unsigned(integer(my_rom(1187)),16);
when x"4a4" => lut_sig <= to_unsigned(integer(my_rom(1188)),16);
when x"4a5" => lut_sig <= to_unsigned(integer(my_rom(1189)),16);
when x"4a6" => lut_sig <= to_unsigned(integer(my_rom(1190)),16);
when x"4a7" => lut_sig <= to_unsigned(integer(my_rom(1191)),16);
when x"4a8" => lut_sig <= to_unsigned(integer(my_rom(1192)),16);
when x"4a9" => lut_sig <= to_unsigned(integer(my_rom(1193)),16);
when x"4aa" => lut_sig <= to_unsigned(integer(my_rom(1194)),16);
when x"4ab" => lut_sig <= to_unsigned(integer(my_rom(1195)),16);
when x"4ac" => lut_sig <= to_unsigned(integer(my_rom(1196)),16);
when x"4ad" => lut_sig <= to_unsigned(integer(my_rom(1197)),16);
when x"4ae" => lut_sig <= to_unsigned(integer(my_rom(1198)),16);
when x"4af" => lut_sig <= to_unsigned(integer(my_rom(1199)),16);
when x"4b0" => lut_sig <= to_unsigned(integer(my_rom(1200)),16);
when x"4b1" => lut_sig <= to_unsigned(integer(my_rom(1201)),16);
when x"4b2" => lut_sig <= to_unsigned(integer(my_rom(1202)),16);
when x"4b3" => lut_sig <= to_unsigned(integer(my_rom(1203)),16);
when x"4b4" => lut_sig <= to_unsigned(integer(my_rom(1204)),16);
when x"4b5" => lut_sig <= to_unsigned(integer(my_rom(1205)),16);
when x"4b6" => lut_sig <= to_unsigned(integer(my_rom(1206)),16);
when x"4b7" => lut_sig <= to_unsigned(integer(my_rom(1207)),16);
when x"4b8" => lut_sig <= to_unsigned(integer(my_rom(1208)),16);
when x"4b9" => lut_sig <= to_unsigned(integer(my_rom(1209)),16);
when x"4ba" => lut_sig <= to_unsigned(integer(my_rom(1210)),16);
when x"4bb" => lut_sig <= to_unsigned(integer(my_rom(1211)),16);
when x"4bc" => lut_sig <= to_unsigned(integer(my_rom(1212)),16);
when x"4bd" => lut_sig <= to_unsigned(integer(my_rom(1213)),16);
when x"4be" => lut_sig <= to_unsigned(integer(my_rom(1214)),16);
when x"4bf" => lut_sig <= to_unsigned(integer(my_rom(1215)),16);
when x"4c0" => lut_sig <= to_unsigned(integer(my_rom(1216)),16);
when x"4c1" => lut_sig <= to_unsigned(integer(my_rom(1217)),16);
when x"4c2" => lut_sig <= to_unsigned(integer(my_rom(1218)),16);
when x"4c3" => lut_sig <= to_unsigned(integer(my_rom(1219)),16);
when x"4c4" => lut_sig <= to_unsigned(integer(my_rom(1220)),16);
when x"4c5" => lut_sig <= to_unsigned(integer(my_rom(1221)),16);
when x"4c6" => lut_sig <= to_unsigned(integer(my_rom(1222)),16);
when x"4c7" => lut_sig <= to_unsigned(integer(my_rom(1223)),16);
when x"4c8" => lut_sig <= to_unsigned(integer(my_rom(1224)),16);
when x"4c9" => lut_sig <= to_unsigned(integer(my_rom(1225)),16);
when x"4ca" => lut_sig <= to_unsigned(integer(my_rom(1226)),16);
when x"4cb" => lut_sig <= to_unsigned(integer(my_rom(1227)),16);
when x"4cc" => lut_sig <= to_unsigned(integer(my_rom(1228)),16);
when x"4cd" => lut_sig <= to_unsigned(integer(my_rom(1229)),16);
when x"4ce" => lut_sig <= to_unsigned(integer(my_rom(1230)),16);
when x"4cf" => lut_sig <= to_unsigned(integer(my_rom(1231)),16);
when x"4d0" => lut_sig <= to_unsigned(integer(my_rom(1232)),16);
when x"4d1" => lut_sig <= to_unsigned(integer(my_rom(1233)),16);
when x"4d2" => lut_sig <= to_unsigned(integer(my_rom(1234)),16);
when x"4d3" => lut_sig <= to_unsigned(integer(my_rom(1235)),16);
when x"4d4" => lut_sig <= to_unsigned(integer(my_rom(1236)),16);
when x"4d5" => lut_sig <= to_unsigned(integer(my_rom(1237)),16);
when x"4d6" => lut_sig <= to_unsigned(integer(my_rom(1238)),16);
when x"4d7" => lut_sig <= to_unsigned(integer(my_rom(1239)),16);
when x"4d8" => lut_sig <= to_unsigned(integer(my_rom(1240)),16);
when x"4d9" => lut_sig <= to_unsigned(integer(my_rom(1241)),16);
when x"4da" => lut_sig <= to_unsigned(integer(my_rom(1242)),16);
when x"4db" => lut_sig <= to_unsigned(integer(my_rom(1243)),16);
when x"4dc" => lut_sig <= to_unsigned(integer(my_rom(1244)),16);
when x"4dd" => lut_sig <= to_unsigned(integer(my_rom(1245)),16);
when x"4de" => lut_sig <= to_unsigned(integer(my_rom(1246)),16);
when x"4df" => lut_sig <= to_unsigned(integer(my_rom(1247)),16);
when x"4e0" => lut_sig <= to_unsigned(integer(my_rom(1248)),16);
when x"4e1" => lut_sig <= to_unsigned(integer(my_rom(1249)),16);
when x"4e2" => lut_sig <= to_unsigned(integer(my_rom(1250)),16);
when x"4e3" => lut_sig <= to_unsigned(integer(my_rom(1251)),16);
when x"4e4" => lut_sig <= to_unsigned(integer(my_rom(1252)),16);
when x"4e5" => lut_sig <= to_unsigned(integer(my_rom(1253)),16);
when x"4e6" => lut_sig <= to_unsigned(integer(my_rom(1254)),16);
when x"4e7" => lut_sig <= to_unsigned(integer(my_rom(1255)),16);
when x"4e8" => lut_sig <= to_unsigned(integer(my_rom(1256)),16);
when x"4e9" => lut_sig <= to_unsigned(integer(my_rom(1257)),16);
when x"4ea" => lut_sig <= to_unsigned(integer(my_rom(1258)),16);
when x"4eb" => lut_sig <= to_unsigned(integer(my_rom(1259)),16);
when x"4ec" => lut_sig <= to_unsigned(integer(my_rom(1260)),16);
when x"4ed" => lut_sig <= to_unsigned(integer(my_rom(1261)),16);
when x"4ee" => lut_sig <= to_unsigned(integer(my_rom(1262)),16);
when x"4ef" => lut_sig <= to_unsigned(integer(my_rom(1263)),16);
when x"4f0" => lut_sig <= to_unsigned(integer(my_rom(1264)),16);
when x"4f1" => lut_sig <= to_unsigned(integer(my_rom(1265)),16);
when x"4f2" => lut_sig <= to_unsigned(integer(my_rom(1266)),16);
when x"4f3" => lut_sig <= to_unsigned(integer(my_rom(1267)),16);
when x"4f4" => lut_sig <= to_unsigned(integer(my_rom(1268)),16);
when x"4f5" => lut_sig <= to_unsigned(integer(my_rom(1269)),16);
when x"4f6" => lut_sig <= to_unsigned(integer(my_rom(1270)),16);
when x"4f7" => lut_sig <= to_unsigned(integer(my_rom(1271)),16);
when x"4f8" => lut_sig <= to_unsigned(integer(my_rom(1272)),16);
when x"4f9" => lut_sig <= to_unsigned(integer(my_rom(1273)),16);
when x"4fa" => lut_sig <= to_unsigned(integer(my_rom(1274)),16);
when x"4fb" => lut_sig <= to_unsigned(integer(my_rom(1275)),16);
when x"4fc" => lut_sig <= to_unsigned(integer(my_rom(1276)),16);
when x"4fd" => lut_sig <= to_unsigned(integer(my_rom(1277)),16);
when x"4fe" => lut_sig <= to_unsigned(integer(my_rom(1278)),16);
when x"4ff" => lut_sig <= to_unsigned(integer(my_rom(1279)),16);
when x"500" => lut_sig <= to_unsigned(integer(my_rom(1280)),16);
when x"501" => lut_sig <= to_unsigned(integer(my_rom(1281)),16);
when x"502" => lut_sig <= to_unsigned(integer(my_rom(1282)),16);
when x"503" => lut_sig <= to_unsigned(integer(my_rom(1283)),16);
when x"504" => lut_sig <= to_unsigned(integer(my_rom(1284)),16);
when x"505" => lut_sig <= to_unsigned(integer(my_rom(1285)),16);
when x"506" => lut_sig <= to_unsigned(integer(my_rom(1286)),16);
when x"507" => lut_sig <= to_unsigned(integer(my_rom(1287)),16);
when x"508" => lut_sig <= to_unsigned(integer(my_rom(1288)),16);
when x"509" => lut_sig <= to_unsigned(integer(my_rom(1289)),16);
when x"50a" => lut_sig <= to_unsigned(integer(my_rom(1290)),16);
when x"50b" => lut_sig <= to_unsigned(integer(my_rom(1291)),16);
when x"50c" => lut_sig <= to_unsigned(integer(my_rom(1292)),16);
when x"50d" => lut_sig <= to_unsigned(integer(my_rom(1293)),16);
when x"50e" => lut_sig <= to_unsigned(integer(my_rom(1294)),16);
when x"50f" => lut_sig <= to_unsigned(integer(my_rom(1295)),16);
when x"510" => lut_sig <= to_unsigned(integer(my_rom(1296)),16);
when x"511" => lut_sig <= to_unsigned(integer(my_rom(1297)),16);
when x"512" => lut_sig <= to_unsigned(integer(my_rom(1298)),16);
when x"513" => lut_sig <= to_unsigned(integer(my_rom(1299)),16);
when x"514" => lut_sig <= to_unsigned(integer(my_rom(1300)),16);
when x"515" => lut_sig <= to_unsigned(integer(my_rom(1301)),16);
when x"516" => lut_sig <= to_unsigned(integer(my_rom(1302)),16);
when x"517" => lut_sig <= to_unsigned(integer(my_rom(1303)),16);
when x"518" => lut_sig <= to_unsigned(integer(my_rom(1304)),16);
when x"519" => lut_sig <= to_unsigned(integer(my_rom(1305)),16);
when x"51a" => lut_sig <= to_unsigned(integer(my_rom(1306)),16);
when x"51b" => lut_sig <= to_unsigned(integer(my_rom(1307)),16);
when x"51c" => lut_sig <= to_unsigned(integer(my_rom(1308)),16);
when x"51d" => lut_sig <= to_unsigned(integer(my_rom(1309)),16);
when x"51e" => lut_sig <= to_unsigned(integer(my_rom(1310)),16);
when x"51f" => lut_sig <= to_unsigned(integer(my_rom(1311)),16);
when x"520" => lut_sig <= to_unsigned(integer(my_rom(1312)),16);
when x"521" => lut_sig <= to_unsigned(integer(my_rom(1313)),16);
when x"522" => lut_sig <= to_unsigned(integer(my_rom(1314)),16);
when x"523" => lut_sig <= to_unsigned(integer(my_rom(1315)),16);
when x"524" => lut_sig <= to_unsigned(integer(my_rom(1316)),16);
when x"525" => lut_sig <= to_unsigned(integer(my_rom(1317)),16);
when x"526" => lut_sig <= to_unsigned(integer(my_rom(1318)),16);
when x"527" => lut_sig <= to_unsigned(integer(my_rom(1319)),16);
when x"528" => lut_sig <= to_unsigned(integer(my_rom(1320)),16);
when x"529" => lut_sig <= to_unsigned(integer(my_rom(1321)),16);
when x"52a" => lut_sig <= to_unsigned(integer(my_rom(1322)),16);
when x"52b" => lut_sig <= to_unsigned(integer(my_rom(1323)),16);
when x"52c" => lut_sig <= to_unsigned(integer(my_rom(1324)),16);
when x"52d" => lut_sig <= to_unsigned(integer(my_rom(1325)),16);
when x"52e" => lut_sig <= to_unsigned(integer(my_rom(1326)),16);
when x"52f" => lut_sig <= to_unsigned(integer(my_rom(1327)),16);
when x"530" => lut_sig <= to_unsigned(integer(my_rom(1328)),16);
when x"531" => lut_sig <= to_unsigned(integer(my_rom(1329)),16);
when x"532" => lut_sig <= to_unsigned(integer(my_rom(1330)),16);
when x"533" => lut_sig <= to_unsigned(integer(my_rom(1331)),16);
when x"534" => lut_sig <= to_unsigned(integer(my_rom(1332)),16);
when x"535" => lut_sig <= to_unsigned(integer(my_rom(1333)),16);
when x"536" => lut_sig <= to_unsigned(integer(my_rom(1334)),16);
when x"537" => lut_sig <= to_unsigned(integer(my_rom(1335)),16);
when x"538" => lut_sig <= to_unsigned(integer(my_rom(1336)),16);
when x"539" => lut_sig <= to_unsigned(integer(my_rom(1337)),16);
when x"53a" => lut_sig <= to_unsigned(integer(my_rom(1338)),16);
when x"53b" => lut_sig <= to_unsigned(integer(my_rom(1339)),16);
when x"53c" => lut_sig <= to_unsigned(integer(my_rom(1340)),16);
when x"53d" => lut_sig <= to_unsigned(integer(my_rom(1341)),16);
when x"53e" => lut_sig <= to_unsigned(integer(my_rom(1342)),16);
when x"53f" => lut_sig <= to_unsigned(integer(my_rom(1343)),16);
when x"540" => lut_sig <= to_unsigned(integer(my_rom(1344)),16);
when x"541" => lut_sig <= to_unsigned(integer(my_rom(1345)),16);
when x"542" => lut_sig <= to_unsigned(integer(my_rom(1346)),16);
when x"543" => lut_sig <= to_unsigned(integer(my_rom(1347)),16);
when x"544" => lut_sig <= to_unsigned(integer(my_rom(1348)),16);
when x"545" => lut_sig <= to_unsigned(integer(my_rom(1349)),16);
when x"546" => lut_sig <= to_unsigned(integer(my_rom(1350)),16);
when x"547" => lut_sig <= to_unsigned(integer(my_rom(1351)),16);
when x"548" => lut_sig <= to_unsigned(integer(my_rom(1352)),16);
when x"549" => lut_sig <= to_unsigned(integer(my_rom(1353)),16);
when x"54a" => lut_sig <= to_unsigned(integer(my_rom(1354)),16);
when x"54b" => lut_sig <= to_unsigned(integer(my_rom(1355)),16);
when x"54c" => lut_sig <= to_unsigned(integer(my_rom(1356)),16);
when x"54d" => lut_sig <= to_unsigned(integer(my_rom(1357)),16);
when x"54e" => lut_sig <= to_unsigned(integer(my_rom(1358)),16);
when x"54f" => lut_sig <= to_unsigned(integer(my_rom(1359)),16);
when x"550" => lut_sig <= to_unsigned(integer(my_rom(1360)),16);
when x"551" => lut_sig <= to_unsigned(integer(my_rom(1361)),16);
when x"552" => lut_sig <= to_unsigned(integer(my_rom(1362)),16);
when x"553" => lut_sig <= to_unsigned(integer(my_rom(1363)),16);
when x"554" => lut_sig <= to_unsigned(integer(my_rom(1364)),16);
when x"555" => lut_sig <= to_unsigned(integer(my_rom(1365)),16);
when x"556" => lut_sig <= to_unsigned(integer(my_rom(1366)),16);
when x"557" => lut_sig <= to_unsigned(integer(my_rom(1367)),16);
when x"558" => lut_sig <= to_unsigned(integer(my_rom(1368)),16);
when x"559" => lut_sig <= to_unsigned(integer(my_rom(1369)),16);
when x"55a" => lut_sig <= to_unsigned(integer(my_rom(1370)),16);
when x"55b" => lut_sig <= to_unsigned(integer(my_rom(1371)),16);
when x"55c" => lut_sig <= to_unsigned(integer(my_rom(1372)),16);
when x"55d" => lut_sig <= to_unsigned(integer(my_rom(1373)),16);
when x"55e" => lut_sig <= to_unsigned(integer(my_rom(1374)),16);
when x"55f" => lut_sig <= to_unsigned(integer(my_rom(1375)),16);
when x"560" => lut_sig <= to_unsigned(integer(my_rom(1376)),16);
when x"561" => lut_sig <= to_unsigned(integer(my_rom(1377)),16);
when x"562" => lut_sig <= to_unsigned(integer(my_rom(1378)),16);
when x"563" => lut_sig <= to_unsigned(integer(my_rom(1379)),16);
when x"564" => lut_sig <= to_unsigned(integer(my_rom(1380)),16);
when x"565" => lut_sig <= to_unsigned(integer(my_rom(1381)),16);
when x"566" => lut_sig <= to_unsigned(integer(my_rom(1382)),16);
when x"567" => lut_sig <= to_unsigned(integer(my_rom(1383)),16);
when x"568" => lut_sig <= to_unsigned(integer(my_rom(1384)),16);
when x"569" => lut_sig <= to_unsigned(integer(my_rom(1385)),16);
when x"56a" => lut_sig <= to_unsigned(integer(my_rom(1386)),16);
when x"56b" => lut_sig <= to_unsigned(integer(my_rom(1387)),16);
when x"56c" => lut_sig <= to_unsigned(integer(my_rom(1388)),16);
when x"56d" => lut_sig <= to_unsigned(integer(my_rom(1389)),16);
when x"56e" => lut_sig <= to_unsigned(integer(my_rom(1390)),16);
when x"56f" => lut_sig <= to_unsigned(integer(my_rom(1391)),16);
when x"570" => lut_sig <= to_unsigned(integer(my_rom(1392)),16);
when x"571" => lut_sig <= to_unsigned(integer(my_rom(1393)),16);
when x"572" => lut_sig <= to_unsigned(integer(my_rom(1394)),16);
when x"573" => lut_sig <= to_unsigned(integer(my_rom(1395)),16);
when x"574" => lut_sig <= to_unsigned(integer(my_rom(1396)),16);
when x"575" => lut_sig <= to_unsigned(integer(my_rom(1397)),16);
when x"576" => lut_sig <= to_unsigned(integer(my_rom(1398)),16);
when x"577" => lut_sig <= to_unsigned(integer(my_rom(1399)),16);
when x"578" => lut_sig <= to_unsigned(integer(my_rom(1400)),16);
when x"579" => lut_sig <= to_unsigned(integer(my_rom(1401)),16);
when x"57a" => lut_sig <= to_unsigned(integer(my_rom(1402)),16);
when x"57b" => lut_sig <= to_unsigned(integer(my_rom(1403)),16);
when x"57c" => lut_sig <= to_unsigned(integer(my_rom(1404)),16);
when x"57d" => lut_sig <= to_unsigned(integer(my_rom(1405)),16);
when x"57e" => lut_sig <= to_unsigned(integer(my_rom(1406)),16);
when x"57f" => lut_sig <= to_unsigned(integer(my_rom(1407)),16);
when x"580" => lut_sig <= to_unsigned(integer(my_rom(1408)),16);
when x"581" => lut_sig <= to_unsigned(integer(my_rom(1409)),16);
when x"582" => lut_sig <= to_unsigned(integer(my_rom(1410)),16);
when x"583" => lut_sig <= to_unsigned(integer(my_rom(1411)),16);
when x"584" => lut_sig <= to_unsigned(integer(my_rom(1412)),16);
when x"585" => lut_sig <= to_unsigned(integer(my_rom(1413)),16);
when x"586" => lut_sig <= to_unsigned(integer(my_rom(1414)),16);
when x"587" => lut_sig <= to_unsigned(integer(my_rom(1415)),16);
when x"588" => lut_sig <= to_unsigned(integer(my_rom(1416)),16);
when x"589" => lut_sig <= to_unsigned(integer(my_rom(1417)),16);
when x"58a" => lut_sig <= to_unsigned(integer(my_rom(1418)),16);
when x"58b" => lut_sig <= to_unsigned(integer(my_rom(1419)),16);
when x"58c" => lut_sig <= to_unsigned(integer(my_rom(1420)),16);
when x"58d" => lut_sig <= to_unsigned(integer(my_rom(1421)),16);
when x"58e" => lut_sig <= to_unsigned(integer(my_rom(1422)),16);
when x"58f" => lut_sig <= to_unsigned(integer(my_rom(1423)),16);
when x"590" => lut_sig <= to_unsigned(integer(my_rom(1424)),16);
when x"591" => lut_sig <= to_unsigned(integer(my_rom(1425)),16);
when x"592" => lut_sig <= to_unsigned(integer(my_rom(1426)),16);
when x"593" => lut_sig <= to_unsigned(integer(my_rom(1427)),16);
when x"594" => lut_sig <= to_unsigned(integer(my_rom(1428)),16);
when x"595" => lut_sig <= to_unsigned(integer(my_rom(1429)),16);
when x"596" => lut_sig <= to_unsigned(integer(my_rom(1430)),16);
when x"597" => lut_sig <= to_unsigned(integer(my_rom(1431)),16);
when x"598" => lut_sig <= to_unsigned(integer(my_rom(1432)),16);
when x"599" => lut_sig <= to_unsigned(integer(my_rom(1433)),16);
when x"59a" => lut_sig <= to_unsigned(integer(my_rom(1434)),16);
when x"59b" => lut_sig <= to_unsigned(integer(my_rom(1435)),16);
when x"59c" => lut_sig <= to_unsigned(integer(my_rom(1436)),16);
when x"59d" => lut_sig <= to_unsigned(integer(my_rom(1437)),16);
when x"59e" => lut_sig <= to_unsigned(integer(my_rom(1438)),16);
when x"59f" => lut_sig <= to_unsigned(integer(my_rom(1439)),16);
when x"5a0" => lut_sig <= to_unsigned(integer(my_rom(1440)),16);
when x"5a1" => lut_sig <= to_unsigned(integer(my_rom(1441)),16);
when x"5a2" => lut_sig <= to_unsigned(integer(my_rom(1442)),16);
when x"5a3" => lut_sig <= to_unsigned(integer(my_rom(1443)),16);
when x"5a4" => lut_sig <= to_unsigned(integer(my_rom(1444)),16);
when x"5a5" => lut_sig <= to_unsigned(integer(my_rom(1445)),16);
when x"5a6" => lut_sig <= to_unsigned(integer(my_rom(1446)),16);
when x"5a7" => lut_sig <= to_unsigned(integer(my_rom(1447)),16);
when x"5a8" => lut_sig <= to_unsigned(integer(my_rom(1448)),16);
when x"5a9" => lut_sig <= to_unsigned(integer(my_rom(1449)),16);
when x"5aa" => lut_sig <= to_unsigned(integer(my_rom(1450)),16);
when x"5ab" => lut_sig <= to_unsigned(integer(my_rom(1451)),16);
when x"5ac" => lut_sig <= to_unsigned(integer(my_rom(1452)),16);
when x"5ad" => lut_sig <= to_unsigned(integer(my_rom(1453)),16);
when x"5ae" => lut_sig <= to_unsigned(integer(my_rom(1454)),16);
when x"5af" => lut_sig <= to_unsigned(integer(my_rom(1455)),16);
when x"5b0" => lut_sig <= to_unsigned(integer(my_rom(1456)),16);
when x"5b1" => lut_sig <= to_unsigned(integer(my_rom(1457)),16);
when x"5b2" => lut_sig <= to_unsigned(integer(my_rom(1458)),16);
when x"5b3" => lut_sig <= to_unsigned(integer(my_rom(1459)),16);
when x"5b4" => lut_sig <= to_unsigned(integer(my_rom(1460)),16);
when x"5b5" => lut_sig <= to_unsigned(integer(my_rom(1461)),16);
when x"5b6" => lut_sig <= to_unsigned(integer(my_rom(1462)),16);
when x"5b7" => lut_sig <= to_unsigned(integer(my_rom(1463)),16);
when x"5b8" => lut_sig <= to_unsigned(integer(my_rom(1464)),16);
when x"5b9" => lut_sig <= to_unsigned(integer(my_rom(1465)),16);
when x"5ba" => lut_sig <= to_unsigned(integer(my_rom(1466)),16);
when x"5bb" => lut_sig <= to_unsigned(integer(my_rom(1467)),16);
when x"5bc" => lut_sig <= to_unsigned(integer(my_rom(1468)),16);
when x"5bd" => lut_sig <= to_unsigned(integer(my_rom(1469)),16);
when x"5be" => lut_sig <= to_unsigned(integer(my_rom(1470)),16);
when x"5bf" => lut_sig <= to_unsigned(integer(my_rom(1471)),16);
when x"5c0" => lut_sig <= to_unsigned(integer(my_rom(1472)),16);
when x"5c1" => lut_sig <= to_unsigned(integer(my_rom(1473)),16);
when x"5c2" => lut_sig <= to_unsigned(integer(my_rom(1474)),16);
when x"5c3" => lut_sig <= to_unsigned(integer(my_rom(1475)),16);
when x"5c4" => lut_sig <= to_unsigned(integer(my_rom(1476)),16);
when x"5c5" => lut_sig <= to_unsigned(integer(my_rom(1477)),16);
when x"5c6" => lut_sig <= to_unsigned(integer(my_rom(1478)),16);
when x"5c7" => lut_sig <= to_unsigned(integer(my_rom(1479)),16);
when x"5c8" => lut_sig <= to_unsigned(integer(my_rom(1480)),16);
when x"5c9" => lut_sig <= to_unsigned(integer(my_rom(1481)),16);
when x"5ca" => lut_sig <= to_unsigned(integer(my_rom(1482)),16);
when x"5cb" => lut_sig <= to_unsigned(integer(my_rom(1483)),16);
when x"5cc" => lut_sig <= to_unsigned(integer(my_rom(1484)),16);
when x"5cd" => lut_sig <= to_unsigned(integer(my_rom(1485)),16);
when x"5ce" => lut_sig <= to_unsigned(integer(my_rom(1486)),16);
when x"5cf" => lut_sig <= to_unsigned(integer(my_rom(1487)),16);
when x"5d0" => lut_sig <= to_unsigned(integer(my_rom(1488)),16);
when x"5d1" => lut_sig <= to_unsigned(integer(my_rom(1489)),16);
when x"5d2" => lut_sig <= to_unsigned(integer(my_rom(1490)),16);
when x"5d3" => lut_sig <= to_unsigned(integer(my_rom(1491)),16);
when x"5d4" => lut_sig <= to_unsigned(integer(my_rom(1492)),16);
when x"5d5" => lut_sig <= to_unsigned(integer(my_rom(1493)),16);
when x"5d6" => lut_sig <= to_unsigned(integer(my_rom(1494)),16);
when x"5d7" => lut_sig <= to_unsigned(integer(my_rom(1495)),16);
when x"5d8" => lut_sig <= to_unsigned(integer(my_rom(1496)),16);
when x"5d9" => lut_sig <= to_unsigned(integer(my_rom(1497)),16);
when x"5da" => lut_sig <= to_unsigned(integer(my_rom(1498)),16);
when x"5db" => lut_sig <= to_unsigned(integer(my_rom(1499)),16);
when x"5dc" => lut_sig <= to_unsigned(integer(my_rom(1500)),16);
when x"5dd" => lut_sig <= to_unsigned(integer(my_rom(1501)),16);
when x"5de" => lut_sig <= to_unsigned(integer(my_rom(1502)),16);
when x"5df" => lut_sig <= to_unsigned(integer(my_rom(1503)),16);
when x"5e0" => lut_sig <= to_unsigned(integer(my_rom(1504)),16);
when x"5e1" => lut_sig <= to_unsigned(integer(my_rom(1505)),16);
when x"5e2" => lut_sig <= to_unsigned(integer(my_rom(1506)),16);
when x"5e3" => lut_sig <= to_unsigned(integer(my_rom(1507)),16);
when x"5e4" => lut_sig <= to_unsigned(integer(my_rom(1508)),16);
when x"5e5" => lut_sig <= to_unsigned(integer(my_rom(1509)),16);
when x"5e6" => lut_sig <= to_unsigned(integer(my_rom(1510)),16);
when x"5e7" => lut_sig <= to_unsigned(integer(my_rom(1511)),16);
when x"5e8" => lut_sig <= to_unsigned(integer(my_rom(1512)),16);
when x"5e9" => lut_sig <= to_unsigned(integer(my_rom(1513)),16);
when x"5ea" => lut_sig <= to_unsigned(integer(my_rom(1514)),16);
when x"5eb" => lut_sig <= to_unsigned(integer(my_rom(1515)),16);
when x"5ec" => lut_sig <= to_unsigned(integer(my_rom(1516)),16);
when x"5ed" => lut_sig <= to_unsigned(integer(my_rom(1517)),16);
when x"5ee" => lut_sig <= to_unsigned(integer(my_rom(1518)),16);
when x"5ef" => lut_sig <= to_unsigned(integer(my_rom(1519)),16);
when x"5f0" => lut_sig <= to_unsigned(integer(my_rom(1520)),16);
when x"5f1" => lut_sig <= to_unsigned(integer(my_rom(1521)),16);
when x"5f2" => lut_sig <= to_unsigned(integer(my_rom(1522)),16);
when x"5f3" => lut_sig <= to_unsigned(integer(my_rom(1523)),16);
when x"5f4" => lut_sig <= to_unsigned(integer(my_rom(1524)),16);
when x"5f5" => lut_sig <= to_unsigned(integer(my_rom(1525)),16);
when x"5f6" => lut_sig <= to_unsigned(integer(my_rom(1526)),16);
when x"5f7" => lut_sig <= to_unsigned(integer(my_rom(1527)),16);
when x"5f8" => lut_sig <= to_unsigned(integer(my_rom(1528)),16);
when x"5f9" => lut_sig <= to_unsigned(integer(my_rom(1529)),16);
when x"5fa" => lut_sig <= to_unsigned(integer(my_rom(1530)),16);
when x"5fb" => lut_sig <= to_unsigned(integer(my_rom(1531)),16);
when x"5fc" => lut_sig <= to_unsigned(integer(my_rom(1532)),16);
when x"5fd" => lut_sig <= to_unsigned(integer(my_rom(1533)),16);
when x"5fe" => lut_sig <= to_unsigned(integer(my_rom(1534)),16);
when x"5ff" => lut_sig <= to_unsigned(integer(my_rom(1535)),16);
when x"600" => lut_sig <= to_unsigned(integer(my_rom(1536)),16);
when x"601" => lut_sig <= to_unsigned(integer(my_rom(1537)),16);
when x"602" => lut_sig <= to_unsigned(integer(my_rom(1538)),16);
when x"603" => lut_sig <= to_unsigned(integer(my_rom(1539)),16);
when x"604" => lut_sig <= to_unsigned(integer(my_rom(1540)),16);
when x"605" => lut_sig <= to_unsigned(integer(my_rom(1541)),16);
when x"606" => lut_sig <= to_unsigned(integer(my_rom(1542)),16);
when x"607" => lut_sig <= to_unsigned(integer(my_rom(1543)),16);
when x"608" => lut_sig <= to_unsigned(integer(my_rom(1544)),16);
when x"609" => lut_sig <= to_unsigned(integer(my_rom(1545)),16);
when x"60a" => lut_sig <= to_unsigned(integer(my_rom(1546)),16);
when x"60b" => lut_sig <= to_unsigned(integer(my_rom(1547)),16);
when x"60c" => lut_sig <= to_unsigned(integer(my_rom(1548)),16);
when x"60d" => lut_sig <= to_unsigned(integer(my_rom(1549)),16);
when x"60e" => lut_sig <= to_unsigned(integer(my_rom(1550)),16);
when x"60f" => lut_sig <= to_unsigned(integer(my_rom(1551)),16);
when x"610" => lut_sig <= to_unsigned(integer(my_rom(1552)),16);
when x"611" => lut_sig <= to_unsigned(integer(my_rom(1553)),16);
when x"612" => lut_sig <= to_unsigned(integer(my_rom(1554)),16);
when x"613" => lut_sig <= to_unsigned(integer(my_rom(1555)),16);
when x"614" => lut_sig <= to_unsigned(integer(my_rom(1556)),16);
when x"615" => lut_sig <= to_unsigned(integer(my_rom(1557)),16);
when x"616" => lut_sig <= to_unsigned(integer(my_rom(1558)),16);
when x"617" => lut_sig <= to_unsigned(integer(my_rom(1559)),16);
when x"618" => lut_sig <= to_unsigned(integer(my_rom(1560)),16);
when x"619" => lut_sig <= to_unsigned(integer(my_rom(1561)),16);
when x"61a" => lut_sig <= to_unsigned(integer(my_rom(1562)),16);
when x"61b" => lut_sig <= to_unsigned(integer(my_rom(1563)),16);
when x"61c" => lut_sig <= to_unsigned(integer(my_rom(1564)),16);
when x"61d" => lut_sig <= to_unsigned(integer(my_rom(1565)),16);
when x"61e" => lut_sig <= to_unsigned(integer(my_rom(1566)),16);
when x"61f" => lut_sig <= to_unsigned(integer(my_rom(1567)),16);
when x"620" => lut_sig <= to_unsigned(integer(my_rom(1568)),16);
when x"621" => lut_sig <= to_unsigned(integer(my_rom(1569)),16);
when x"622" => lut_sig <= to_unsigned(integer(my_rom(1570)),16);
when x"623" => lut_sig <= to_unsigned(integer(my_rom(1571)),16);
when x"624" => lut_sig <= to_unsigned(integer(my_rom(1572)),16);
when x"625" => lut_sig <= to_unsigned(integer(my_rom(1573)),16);
when x"626" => lut_sig <= to_unsigned(integer(my_rom(1574)),16);
when x"627" => lut_sig <= to_unsigned(integer(my_rom(1575)),16);
when x"628" => lut_sig <= to_unsigned(integer(my_rom(1576)),16);
when x"629" => lut_sig <= to_unsigned(integer(my_rom(1577)),16);
when x"62a" => lut_sig <= to_unsigned(integer(my_rom(1578)),16);
when x"62b" => lut_sig <= to_unsigned(integer(my_rom(1579)),16);
when x"62c" => lut_sig <= to_unsigned(integer(my_rom(1580)),16);
when x"62d" => lut_sig <= to_unsigned(integer(my_rom(1581)),16);
when x"62e" => lut_sig <= to_unsigned(integer(my_rom(1582)),16);
when x"62f" => lut_sig <= to_unsigned(integer(my_rom(1583)),16);
when x"630" => lut_sig <= to_unsigned(integer(my_rom(1584)),16);
when x"631" => lut_sig <= to_unsigned(integer(my_rom(1585)),16);
when x"632" => lut_sig <= to_unsigned(integer(my_rom(1586)),16);
when x"633" => lut_sig <= to_unsigned(integer(my_rom(1587)),16);
when x"634" => lut_sig <= to_unsigned(integer(my_rom(1588)),16);
when x"635" => lut_sig <= to_unsigned(integer(my_rom(1589)),16);
when x"636" => lut_sig <= to_unsigned(integer(my_rom(1590)),16);
when x"637" => lut_sig <= to_unsigned(integer(my_rom(1591)),16);
when x"638" => lut_sig <= to_unsigned(integer(my_rom(1592)),16);
when x"639" => lut_sig <= to_unsigned(integer(my_rom(1593)),16);
when x"63a" => lut_sig <= to_unsigned(integer(my_rom(1594)),16);
when x"63b" => lut_sig <= to_unsigned(integer(my_rom(1595)),16);
when x"63c" => lut_sig <= to_unsigned(integer(my_rom(1596)),16);
when x"63d" => lut_sig <= to_unsigned(integer(my_rom(1597)),16);
when x"63e" => lut_sig <= to_unsigned(integer(my_rom(1598)),16);
when x"63f" => lut_sig <= to_unsigned(integer(my_rom(1599)),16);
when x"640" => lut_sig <= to_unsigned(integer(my_rom(1600)),16);
when x"641" => lut_sig <= to_unsigned(integer(my_rom(1601)),16);
when x"642" => lut_sig <= to_unsigned(integer(my_rom(1602)),16);
when x"643" => lut_sig <= to_unsigned(integer(my_rom(1603)),16);
when x"644" => lut_sig <= to_unsigned(integer(my_rom(1604)),16);
when x"645" => lut_sig <= to_unsigned(integer(my_rom(1605)),16);
when x"646" => lut_sig <= to_unsigned(integer(my_rom(1606)),16);
when x"647" => lut_sig <= to_unsigned(integer(my_rom(1607)),16);
when x"648" => lut_sig <= to_unsigned(integer(my_rom(1608)),16);
when x"649" => lut_sig <= to_unsigned(integer(my_rom(1609)),16);
when x"64a" => lut_sig <= to_unsigned(integer(my_rom(1610)),16);
when x"64b" => lut_sig <= to_unsigned(integer(my_rom(1611)),16);
when x"64c" => lut_sig <= to_unsigned(integer(my_rom(1612)),16);
when x"64d" => lut_sig <= to_unsigned(integer(my_rom(1613)),16);
when x"64e" => lut_sig <= to_unsigned(integer(my_rom(1614)),16);
when x"64f" => lut_sig <= to_unsigned(integer(my_rom(1615)),16);
when x"650" => lut_sig <= to_unsigned(integer(my_rom(1616)),16);
when x"651" => lut_sig <= to_unsigned(integer(my_rom(1617)),16);
when x"652" => lut_sig <= to_unsigned(integer(my_rom(1618)),16);
when x"653" => lut_sig <= to_unsigned(integer(my_rom(1619)),16);
when x"654" => lut_sig <= to_unsigned(integer(my_rom(1620)),16);
when x"655" => lut_sig <= to_unsigned(integer(my_rom(1621)),16);
when x"656" => lut_sig <= to_unsigned(integer(my_rom(1622)),16);
when x"657" => lut_sig <= to_unsigned(integer(my_rom(1623)),16);
when x"658" => lut_sig <= to_unsigned(integer(my_rom(1624)),16);
when x"659" => lut_sig <= to_unsigned(integer(my_rom(1625)),16);
when x"65a" => lut_sig <= to_unsigned(integer(my_rom(1626)),16);
when x"65b" => lut_sig <= to_unsigned(integer(my_rom(1627)),16);
when x"65c" => lut_sig <= to_unsigned(integer(my_rom(1628)),16);
when x"65d" => lut_sig <= to_unsigned(integer(my_rom(1629)),16);
when x"65e" => lut_sig <= to_unsigned(integer(my_rom(1630)),16);
when x"65f" => lut_sig <= to_unsigned(integer(my_rom(1631)),16);
when x"660" => lut_sig <= to_unsigned(integer(my_rom(1632)),16);
when x"661" => lut_sig <= to_unsigned(integer(my_rom(1633)),16);
when x"662" => lut_sig <= to_unsigned(integer(my_rom(1634)),16);
when x"663" => lut_sig <= to_unsigned(integer(my_rom(1635)),16);
when x"664" => lut_sig <= to_unsigned(integer(my_rom(1636)),16);
when x"665" => lut_sig <= to_unsigned(integer(my_rom(1637)),16);
when x"666" => lut_sig <= to_unsigned(integer(my_rom(1638)),16);
when x"667" => lut_sig <= to_unsigned(integer(my_rom(1639)),16);
when x"668" => lut_sig <= to_unsigned(integer(my_rom(1640)),16);
when x"669" => lut_sig <= to_unsigned(integer(my_rom(1641)),16);
when x"66a" => lut_sig <= to_unsigned(integer(my_rom(1642)),16);
when x"66b" => lut_sig <= to_unsigned(integer(my_rom(1643)),16);
when x"66c" => lut_sig <= to_unsigned(integer(my_rom(1644)),16);
when x"66d" => lut_sig <= to_unsigned(integer(my_rom(1645)),16);
when x"66e" => lut_sig <= to_unsigned(integer(my_rom(1646)),16);
when x"66f" => lut_sig <= to_unsigned(integer(my_rom(1647)),16);
when x"670" => lut_sig <= to_unsigned(integer(my_rom(1648)),16);
when x"671" => lut_sig <= to_unsigned(integer(my_rom(1649)),16);
when x"672" => lut_sig <= to_unsigned(integer(my_rom(1650)),16);
when x"673" => lut_sig <= to_unsigned(integer(my_rom(1651)),16);
when x"674" => lut_sig <= to_unsigned(integer(my_rom(1652)),16);
when x"675" => lut_sig <= to_unsigned(integer(my_rom(1653)),16);
when x"676" => lut_sig <= to_unsigned(integer(my_rom(1654)),16);
when x"677" => lut_sig <= to_unsigned(integer(my_rom(1655)),16);
when x"678" => lut_sig <= to_unsigned(integer(my_rom(1656)),16);
when x"679" => lut_sig <= to_unsigned(integer(my_rom(1657)),16);
when x"67a" => lut_sig <= to_unsigned(integer(my_rom(1658)),16);
when x"67b" => lut_sig <= to_unsigned(integer(my_rom(1659)),16);
when x"67c" => lut_sig <= to_unsigned(integer(my_rom(1660)),16);
when x"67d" => lut_sig <= to_unsigned(integer(my_rom(1661)),16);
when x"67e" => lut_sig <= to_unsigned(integer(my_rom(1662)),16);
when x"67f" => lut_sig <= to_unsigned(integer(my_rom(1663)),16);
when x"680" => lut_sig <= to_unsigned(integer(my_rom(1664)),16);
when x"681" => lut_sig <= to_unsigned(integer(my_rom(1665)),16);
when x"682" => lut_sig <= to_unsigned(integer(my_rom(1666)),16);
when x"683" => lut_sig <= to_unsigned(integer(my_rom(1667)),16);
when x"684" => lut_sig <= to_unsigned(integer(my_rom(1668)),16);
when x"685" => lut_sig <= to_unsigned(integer(my_rom(1669)),16);
when x"686" => lut_sig <= to_unsigned(integer(my_rom(1670)),16);
when x"687" => lut_sig <= to_unsigned(integer(my_rom(1671)),16);
when x"688" => lut_sig <= to_unsigned(integer(my_rom(1672)),16);
when x"689" => lut_sig <= to_unsigned(integer(my_rom(1673)),16);
when x"68a" => lut_sig <= to_unsigned(integer(my_rom(1674)),16);
when x"68b" => lut_sig <= to_unsigned(integer(my_rom(1675)),16);
when x"68c" => lut_sig <= to_unsigned(integer(my_rom(1676)),16);
when x"68d" => lut_sig <= to_unsigned(integer(my_rom(1677)),16);
when x"68e" => lut_sig <= to_unsigned(integer(my_rom(1678)),16);
when x"68f" => lut_sig <= to_unsigned(integer(my_rom(1679)),16);
when x"690" => lut_sig <= to_unsigned(integer(my_rom(1680)),16);
when x"691" => lut_sig <= to_unsigned(integer(my_rom(1681)),16);
when x"692" => lut_sig <= to_unsigned(integer(my_rom(1682)),16);
when x"693" => lut_sig <= to_unsigned(integer(my_rom(1683)),16);
when x"694" => lut_sig <= to_unsigned(integer(my_rom(1684)),16);
when x"695" => lut_sig <= to_unsigned(integer(my_rom(1685)),16);
when x"696" => lut_sig <= to_unsigned(integer(my_rom(1686)),16);
when x"697" => lut_sig <= to_unsigned(integer(my_rom(1687)),16);
when x"698" => lut_sig <= to_unsigned(integer(my_rom(1688)),16);
when x"699" => lut_sig <= to_unsigned(integer(my_rom(1689)),16);
when x"69a" => lut_sig <= to_unsigned(integer(my_rom(1690)),16);
when x"69b" => lut_sig <= to_unsigned(integer(my_rom(1691)),16);
when x"69c" => lut_sig <= to_unsigned(integer(my_rom(1692)),16);
when x"69d" => lut_sig <= to_unsigned(integer(my_rom(1693)),16);
when x"69e" => lut_sig <= to_unsigned(integer(my_rom(1694)),16);
when x"69f" => lut_sig <= to_unsigned(integer(my_rom(1695)),16);
when x"6a0" => lut_sig <= to_unsigned(integer(my_rom(1696)),16);
when x"6a1" => lut_sig <= to_unsigned(integer(my_rom(1697)),16);
when x"6a2" => lut_sig <= to_unsigned(integer(my_rom(1698)),16);
when x"6a3" => lut_sig <= to_unsigned(integer(my_rom(1699)),16);
when x"6a4" => lut_sig <= to_unsigned(integer(my_rom(1700)),16);
when x"6a5" => lut_sig <= to_unsigned(integer(my_rom(1701)),16);
when x"6a6" => lut_sig <= to_unsigned(integer(my_rom(1702)),16);
when x"6a7" => lut_sig <= to_unsigned(integer(my_rom(1703)),16);
when x"6a8" => lut_sig <= to_unsigned(integer(my_rom(1704)),16);
when x"6a9" => lut_sig <= to_unsigned(integer(my_rom(1705)),16);
when x"6aa" => lut_sig <= to_unsigned(integer(my_rom(1706)),16);
when x"6ab" => lut_sig <= to_unsigned(integer(my_rom(1707)),16);
when x"6ac" => lut_sig <= to_unsigned(integer(my_rom(1708)),16);
when x"6ad" => lut_sig <= to_unsigned(integer(my_rom(1709)),16);
when x"6ae" => lut_sig <= to_unsigned(integer(my_rom(1710)),16);
when x"6af" => lut_sig <= to_unsigned(integer(my_rom(1711)),16);
when x"6b0" => lut_sig <= to_unsigned(integer(my_rom(1712)),16);
when x"6b1" => lut_sig <= to_unsigned(integer(my_rom(1713)),16);
when x"6b2" => lut_sig <= to_unsigned(integer(my_rom(1714)),16);
when x"6b3" => lut_sig <= to_unsigned(integer(my_rom(1715)),16);
when x"6b4" => lut_sig <= to_unsigned(integer(my_rom(1716)),16);
when x"6b5" => lut_sig <= to_unsigned(integer(my_rom(1717)),16);
when x"6b6" => lut_sig <= to_unsigned(integer(my_rom(1718)),16);
when x"6b7" => lut_sig <= to_unsigned(integer(my_rom(1719)),16);
when x"6b8" => lut_sig <= to_unsigned(integer(my_rom(1720)),16);
when x"6b9" => lut_sig <= to_unsigned(integer(my_rom(1721)),16);
when x"6ba" => lut_sig <= to_unsigned(integer(my_rom(1722)),16);
when x"6bb" => lut_sig <= to_unsigned(integer(my_rom(1723)),16);
when x"6bc" => lut_sig <= to_unsigned(integer(my_rom(1724)),16);
when x"6bd" => lut_sig <= to_unsigned(integer(my_rom(1725)),16);
when x"6be" => lut_sig <= to_unsigned(integer(my_rom(1726)),16);
when x"6bf" => lut_sig <= to_unsigned(integer(my_rom(1727)),16);
when x"6c0" => lut_sig <= to_unsigned(integer(my_rom(1728)),16);
when x"6c1" => lut_sig <= to_unsigned(integer(my_rom(1729)),16);
when x"6c2" => lut_sig <= to_unsigned(integer(my_rom(1730)),16);
when x"6c3" => lut_sig <= to_unsigned(integer(my_rom(1731)),16);
when x"6c4" => lut_sig <= to_unsigned(integer(my_rom(1732)),16);
when x"6c5" => lut_sig <= to_unsigned(integer(my_rom(1733)),16);
when x"6c6" => lut_sig <= to_unsigned(integer(my_rom(1734)),16);
when x"6c7" => lut_sig <= to_unsigned(integer(my_rom(1735)),16);
when x"6c8" => lut_sig <= to_unsigned(integer(my_rom(1736)),16);
when x"6c9" => lut_sig <= to_unsigned(integer(my_rom(1737)),16);
when x"6ca" => lut_sig <= to_unsigned(integer(my_rom(1738)),16);
when x"6cb" => lut_sig <= to_unsigned(integer(my_rom(1739)),16);
when x"6cc" => lut_sig <= to_unsigned(integer(my_rom(1740)),16);
when x"6cd" => lut_sig <= to_unsigned(integer(my_rom(1741)),16);
when x"6ce" => lut_sig <= to_unsigned(integer(my_rom(1742)),16);
when x"6cf" => lut_sig <= to_unsigned(integer(my_rom(1743)),16);
when x"6d0" => lut_sig <= to_unsigned(integer(my_rom(1744)),16);
when x"6d1" => lut_sig <= to_unsigned(integer(my_rom(1745)),16);
when x"6d2" => lut_sig <= to_unsigned(integer(my_rom(1746)),16);
when x"6d3" => lut_sig <= to_unsigned(integer(my_rom(1747)),16);
when x"6d4" => lut_sig <= to_unsigned(integer(my_rom(1748)),16);
when x"6d5" => lut_sig <= to_unsigned(integer(my_rom(1749)),16);
when x"6d6" => lut_sig <= to_unsigned(integer(my_rom(1750)),16);
when x"6d7" => lut_sig <= to_unsigned(integer(my_rom(1751)),16);
when x"6d8" => lut_sig <= to_unsigned(integer(my_rom(1752)),16);
when x"6d9" => lut_sig <= to_unsigned(integer(my_rom(1753)),16);
when x"6da" => lut_sig <= to_unsigned(integer(my_rom(1754)),16);
when x"6db" => lut_sig <= to_unsigned(integer(my_rom(1755)),16);
when x"6dc" => lut_sig <= to_unsigned(integer(my_rom(1756)),16);
when x"6dd" => lut_sig <= to_unsigned(integer(my_rom(1757)),16);
when x"6de" => lut_sig <= to_unsigned(integer(my_rom(1758)),16);
when x"6df" => lut_sig <= to_unsigned(integer(my_rom(1759)),16);
when x"6e0" => lut_sig <= to_unsigned(integer(my_rom(1760)),16);
when x"6e1" => lut_sig <= to_unsigned(integer(my_rom(1761)),16);
when x"6e2" => lut_sig <= to_unsigned(integer(my_rom(1762)),16);
when x"6e3" => lut_sig <= to_unsigned(integer(my_rom(1763)),16);
when x"6e4" => lut_sig <= to_unsigned(integer(my_rom(1764)),16);
when x"6e5" => lut_sig <= to_unsigned(integer(my_rom(1765)),16);
when x"6e6" => lut_sig <= to_unsigned(integer(my_rom(1766)),16);
when x"6e7" => lut_sig <= to_unsigned(integer(my_rom(1767)),16);
when x"6e8" => lut_sig <= to_unsigned(integer(my_rom(1768)),16);
when x"6e9" => lut_sig <= to_unsigned(integer(my_rom(1769)),16);
when x"6ea" => lut_sig <= to_unsigned(integer(my_rom(1770)),16);
when x"6eb" => lut_sig <= to_unsigned(integer(my_rom(1771)),16);
when x"6ec" => lut_sig <= to_unsigned(integer(my_rom(1772)),16);
when x"6ed" => lut_sig <= to_unsigned(integer(my_rom(1773)),16);
when x"6ee" => lut_sig <= to_unsigned(integer(my_rom(1774)),16);
when x"6ef" => lut_sig <= to_unsigned(integer(my_rom(1775)),16);
when x"6f0" => lut_sig <= to_unsigned(integer(my_rom(1776)),16);
when x"6f1" => lut_sig <= to_unsigned(integer(my_rom(1777)),16);
when x"6f2" => lut_sig <= to_unsigned(integer(my_rom(1778)),16);
when x"6f3" => lut_sig <= to_unsigned(integer(my_rom(1779)),16);
when x"6f4" => lut_sig <= to_unsigned(integer(my_rom(1780)),16);
when x"6f5" => lut_sig <= to_unsigned(integer(my_rom(1781)),16);
when x"6f6" => lut_sig <= to_unsigned(integer(my_rom(1782)),16);
when x"6f7" => lut_sig <= to_unsigned(integer(my_rom(1783)),16);
when x"6f8" => lut_sig <= to_unsigned(integer(my_rom(1784)),16);
when x"6f9" => lut_sig <= to_unsigned(integer(my_rom(1785)),16);
when x"6fa" => lut_sig <= to_unsigned(integer(my_rom(1786)),16);
when x"6fb" => lut_sig <= to_unsigned(integer(my_rom(1787)),16);
when x"6fc" => lut_sig <= to_unsigned(integer(my_rom(1788)),16);
when x"6fd" => lut_sig <= to_unsigned(integer(my_rom(1789)),16);
when x"6fe" => lut_sig <= to_unsigned(integer(my_rom(1790)),16);
when x"6ff" => lut_sig <= to_unsigned(integer(my_rom(1791)),16);
when x"700" => lut_sig <= to_unsigned(integer(my_rom(1792)),16);
when x"701" => lut_sig <= to_unsigned(integer(my_rom(1793)),16);
when x"702" => lut_sig <= to_unsigned(integer(my_rom(1794)),16);
when x"703" => lut_sig <= to_unsigned(integer(my_rom(1795)),16);
when x"704" => lut_sig <= to_unsigned(integer(my_rom(1796)),16);
when x"705" => lut_sig <= to_unsigned(integer(my_rom(1797)),16);
when x"706" => lut_sig <= to_unsigned(integer(my_rom(1798)),16);
when x"707" => lut_sig <= to_unsigned(integer(my_rom(1799)),16);
when x"708" => lut_sig <= to_unsigned(integer(my_rom(1800)),16);
when x"709" => lut_sig <= to_unsigned(integer(my_rom(1801)),16);
when x"70a" => lut_sig <= to_unsigned(integer(my_rom(1802)),16);
when x"70b" => lut_sig <= to_unsigned(integer(my_rom(1803)),16);
when x"70c" => lut_sig <= to_unsigned(integer(my_rom(1804)),16);
when x"70d" => lut_sig <= to_unsigned(integer(my_rom(1805)),16);
when x"70e" => lut_sig <= to_unsigned(integer(my_rom(1806)),16);
when x"70f" => lut_sig <= to_unsigned(integer(my_rom(1807)),16);
when x"710" => lut_sig <= to_unsigned(integer(my_rom(1808)),16);
when x"711" => lut_sig <= to_unsigned(integer(my_rom(1809)),16);
when x"712" => lut_sig <= to_unsigned(integer(my_rom(1810)),16);
when x"713" => lut_sig <= to_unsigned(integer(my_rom(1811)),16);
when x"714" => lut_sig <= to_unsigned(integer(my_rom(1812)),16);
when x"715" => lut_sig <= to_unsigned(integer(my_rom(1813)),16);
when x"716" => lut_sig <= to_unsigned(integer(my_rom(1814)),16);
when x"717" => lut_sig <= to_unsigned(integer(my_rom(1815)),16);
when x"718" => lut_sig <= to_unsigned(integer(my_rom(1816)),16);
when x"719" => lut_sig <= to_unsigned(integer(my_rom(1817)),16);
when x"71a" => lut_sig <= to_unsigned(integer(my_rom(1818)),16);
when x"71b" => lut_sig <= to_unsigned(integer(my_rom(1819)),16);
when x"71c" => lut_sig <= to_unsigned(integer(my_rom(1820)),16);
when x"71d" => lut_sig <= to_unsigned(integer(my_rom(1821)),16);
when x"71e" => lut_sig <= to_unsigned(integer(my_rom(1822)),16);
when x"71f" => lut_sig <= to_unsigned(integer(my_rom(1823)),16);
when x"720" => lut_sig <= to_unsigned(integer(my_rom(1824)),16);
when x"721" => lut_sig <= to_unsigned(integer(my_rom(1825)),16);
when x"722" => lut_sig <= to_unsigned(integer(my_rom(1826)),16);
when x"723" => lut_sig <= to_unsigned(integer(my_rom(1827)),16);
when x"724" => lut_sig <= to_unsigned(integer(my_rom(1828)),16);
when x"725" => lut_sig <= to_unsigned(integer(my_rom(1829)),16);
when x"726" => lut_sig <= to_unsigned(integer(my_rom(1830)),16);
when x"727" => lut_sig <= to_unsigned(integer(my_rom(1831)),16);
when x"728" => lut_sig <= to_unsigned(integer(my_rom(1832)),16);
when x"729" => lut_sig <= to_unsigned(integer(my_rom(1833)),16);
when x"72a" => lut_sig <= to_unsigned(integer(my_rom(1834)),16);
when x"72b" => lut_sig <= to_unsigned(integer(my_rom(1835)),16);
when x"72c" => lut_sig <= to_unsigned(integer(my_rom(1836)),16);
when x"72d" => lut_sig <= to_unsigned(integer(my_rom(1837)),16);
when x"72e" => lut_sig <= to_unsigned(integer(my_rom(1838)),16);
when x"72f" => lut_sig <= to_unsigned(integer(my_rom(1839)),16);
when x"730" => lut_sig <= to_unsigned(integer(my_rom(1840)),16);
when x"731" => lut_sig <= to_unsigned(integer(my_rom(1841)),16);
when x"732" => lut_sig <= to_unsigned(integer(my_rom(1842)),16);
when x"733" => lut_sig <= to_unsigned(integer(my_rom(1843)),16);
when x"734" => lut_sig <= to_unsigned(integer(my_rom(1844)),16);
when x"735" => lut_sig <= to_unsigned(integer(my_rom(1845)),16);
when x"736" => lut_sig <= to_unsigned(integer(my_rom(1846)),16);
when x"737" => lut_sig <= to_unsigned(integer(my_rom(1847)),16);
when x"738" => lut_sig <= to_unsigned(integer(my_rom(1848)),16);
when x"739" => lut_sig <= to_unsigned(integer(my_rom(1849)),16);
when x"73a" => lut_sig <= to_unsigned(integer(my_rom(1850)),16);
when x"73b" => lut_sig <= to_unsigned(integer(my_rom(1851)),16);
when x"73c" => lut_sig <= to_unsigned(integer(my_rom(1852)),16);
when x"73d" => lut_sig <= to_unsigned(integer(my_rom(1853)),16);
when x"73e" => lut_sig <= to_unsigned(integer(my_rom(1854)),16);
when x"73f" => lut_sig <= to_unsigned(integer(my_rom(1855)),16);
when x"740" => lut_sig <= to_unsigned(integer(my_rom(1856)),16);
when x"741" => lut_sig <= to_unsigned(integer(my_rom(1857)),16);
when x"742" => lut_sig <= to_unsigned(integer(my_rom(1858)),16);
when x"743" => lut_sig <= to_unsigned(integer(my_rom(1859)),16);
when x"744" => lut_sig <= to_unsigned(integer(my_rom(1860)),16);
when x"745" => lut_sig <= to_unsigned(integer(my_rom(1861)),16);
when x"746" => lut_sig <= to_unsigned(integer(my_rom(1862)),16);
when x"747" => lut_sig <= to_unsigned(integer(my_rom(1863)),16);
when x"748" => lut_sig <= to_unsigned(integer(my_rom(1864)),16);
when x"749" => lut_sig <= to_unsigned(integer(my_rom(1865)),16);
when x"74a" => lut_sig <= to_unsigned(integer(my_rom(1866)),16);
when x"74b" => lut_sig <= to_unsigned(integer(my_rom(1867)),16);
when x"74c" => lut_sig <= to_unsigned(integer(my_rom(1868)),16);
when x"74d" => lut_sig <= to_unsigned(integer(my_rom(1869)),16);
when x"74e" => lut_sig <= to_unsigned(integer(my_rom(1870)),16);
when x"74f" => lut_sig <= to_unsigned(integer(my_rom(1871)),16);
when x"750" => lut_sig <= to_unsigned(integer(my_rom(1872)),16);
when x"751" => lut_sig <= to_unsigned(integer(my_rom(1873)),16);
when x"752" => lut_sig <= to_unsigned(integer(my_rom(1874)),16);
when x"753" => lut_sig <= to_unsigned(integer(my_rom(1875)),16);
when x"754" => lut_sig <= to_unsigned(integer(my_rom(1876)),16);
when x"755" => lut_sig <= to_unsigned(integer(my_rom(1877)),16);
when x"756" => lut_sig <= to_unsigned(integer(my_rom(1878)),16);
when x"757" => lut_sig <= to_unsigned(integer(my_rom(1879)),16);
when x"758" => lut_sig <= to_unsigned(integer(my_rom(1880)),16);
when x"759" => lut_sig <= to_unsigned(integer(my_rom(1881)),16);
when x"75a" => lut_sig <= to_unsigned(integer(my_rom(1882)),16);
when x"75b" => lut_sig <= to_unsigned(integer(my_rom(1883)),16);
when x"75c" => lut_sig <= to_unsigned(integer(my_rom(1884)),16);
when x"75d" => lut_sig <= to_unsigned(integer(my_rom(1885)),16);
when x"75e" => lut_sig <= to_unsigned(integer(my_rom(1886)),16);
when x"75f" => lut_sig <= to_unsigned(integer(my_rom(1887)),16);
when x"760" => lut_sig <= to_unsigned(integer(my_rom(1888)),16);
when x"761" => lut_sig <= to_unsigned(integer(my_rom(1889)),16);
when x"762" => lut_sig <= to_unsigned(integer(my_rom(1890)),16);
when x"763" => lut_sig <= to_unsigned(integer(my_rom(1891)),16);
when x"764" => lut_sig <= to_unsigned(integer(my_rom(1892)),16);
when x"765" => lut_sig <= to_unsigned(integer(my_rom(1893)),16);
when x"766" => lut_sig <= to_unsigned(integer(my_rom(1894)),16);
when x"767" => lut_sig <= to_unsigned(integer(my_rom(1895)),16);
when x"768" => lut_sig <= to_unsigned(integer(my_rom(1896)),16);
when x"769" => lut_sig <= to_unsigned(integer(my_rom(1897)),16);
when x"76a" => lut_sig <= to_unsigned(integer(my_rom(1898)),16);
when x"76b" => lut_sig <= to_unsigned(integer(my_rom(1899)),16);
when x"76c" => lut_sig <= to_unsigned(integer(my_rom(1900)),16);
when x"76d" => lut_sig <= to_unsigned(integer(my_rom(1901)),16);
when x"76e" => lut_sig <= to_unsigned(integer(my_rom(1902)),16);
when x"76f" => lut_sig <= to_unsigned(integer(my_rom(1903)),16);
when x"770" => lut_sig <= to_unsigned(integer(my_rom(1904)),16);
when x"771" => lut_sig <= to_unsigned(integer(my_rom(1905)),16);
when x"772" => lut_sig <= to_unsigned(integer(my_rom(1906)),16);
when x"773" => lut_sig <= to_unsigned(integer(my_rom(1907)),16);
when x"774" => lut_sig <= to_unsigned(integer(my_rom(1908)),16);
when x"775" => lut_sig <= to_unsigned(integer(my_rom(1909)),16);
when x"776" => lut_sig <= to_unsigned(integer(my_rom(1910)),16);
when x"777" => lut_sig <= to_unsigned(integer(my_rom(1911)),16);
when x"778" => lut_sig <= to_unsigned(integer(my_rom(1912)),16);
when x"779" => lut_sig <= to_unsigned(integer(my_rom(1913)),16);
when x"77a" => lut_sig <= to_unsigned(integer(my_rom(1914)),16);
when x"77b" => lut_sig <= to_unsigned(integer(my_rom(1915)),16);
when x"77c" => lut_sig <= to_unsigned(integer(my_rom(1916)),16);
when x"77d" => lut_sig <= to_unsigned(integer(my_rom(1917)),16);
when x"77e" => lut_sig <= to_unsigned(integer(my_rom(1918)),16);
when x"77f" => lut_sig <= to_unsigned(integer(my_rom(1919)),16);
when x"780" => lut_sig <= to_unsigned(integer(my_rom(1920)),16);
when x"781" => lut_sig <= to_unsigned(integer(my_rom(1921)),16);
when x"782" => lut_sig <= to_unsigned(integer(my_rom(1922)),16);
when x"783" => lut_sig <= to_unsigned(integer(my_rom(1923)),16);
when x"784" => lut_sig <= to_unsigned(integer(my_rom(1924)),16);
when x"785" => lut_sig <= to_unsigned(integer(my_rom(1925)),16);
when x"786" => lut_sig <= to_unsigned(integer(my_rom(1926)),16);
when x"787" => lut_sig <= to_unsigned(integer(my_rom(1927)),16);
when x"788" => lut_sig <= to_unsigned(integer(my_rom(1928)),16);
when x"789" => lut_sig <= to_unsigned(integer(my_rom(1929)),16);
when x"78a" => lut_sig <= to_unsigned(integer(my_rom(1930)),16);
when x"78b" => lut_sig <= to_unsigned(integer(my_rom(1931)),16);
when x"78c" => lut_sig <= to_unsigned(integer(my_rom(1932)),16);
when x"78d" => lut_sig <= to_unsigned(integer(my_rom(1933)),16);
when x"78e" => lut_sig <= to_unsigned(integer(my_rom(1934)),16);
when x"78f" => lut_sig <= to_unsigned(integer(my_rom(1935)),16);
when x"790" => lut_sig <= to_unsigned(integer(my_rom(1936)),16);
when x"791" => lut_sig <= to_unsigned(integer(my_rom(1937)),16);
when x"792" => lut_sig <= to_unsigned(integer(my_rom(1938)),16);
when x"793" => lut_sig <= to_unsigned(integer(my_rom(1939)),16);
when x"794" => lut_sig <= to_unsigned(integer(my_rom(1940)),16);
when x"795" => lut_sig <= to_unsigned(integer(my_rom(1941)),16);
when x"796" => lut_sig <= to_unsigned(integer(my_rom(1942)),16);
when x"797" => lut_sig <= to_unsigned(integer(my_rom(1943)),16);
when x"798" => lut_sig <= to_unsigned(integer(my_rom(1944)),16);
when x"799" => lut_sig <= to_unsigned(integer(my_rom(1945)),16);
when x"79a" => lut_sig <= to_unsigned(integer(my_rom(1946)),16);
when x"79b" => lut_sig <= to_unsigned(integer(my_rom(1947)),16);
when x"79c" => lut_sig <= to_unsigned(integer(my_rom(1948)),16);
when x"79d" => lut_sig <= to_unsigned(integer(my_rom(1949)),16);
when x"79e" => lut_sig <= to_unsigned(integer(my_rom(1950)),16);
when x"79f" => lut_sig <= to_unsigned(integer(my_rom(1951)),16);
when x"7a0" => lut_sig <= to_unsigned(integer(my_rom(1952)),16);
when x"7a1" => lut_sig <= to_unsigned(integer(my_rom(1953)),16);
when x"7a2" => lut_sig <= to_unsigned(integer(my_rom(1954)),16);
when x"7a3" => lut_sig <= to_unsigned(integer(my_rom(1955)),16);
when x"7a4" => lut_sig <= to_unsigned(integer(my_rom(1956)),16);
when x"7a5" => lut_sig <= to_unsigned(integer(my_rom(1957)),16);
when x"7a6" => lut_sig <= to_unsigned(integer(my_rom(1958)),16);
when x"7a7" => lut_sig <= to_unsigned(integer(my_rom(1959)),16);
when x"7a8" => lut_sig <= to_unsigned(integer(my_rom(1960)),16);
when x"7a9" => lut_sig <= to_unsigned(integer(my_rom(1961)),16);
when x"7aa" => lut_sig <= to_unsigned(integer(my_rom(1962)),16);
when x"7ab" => lut_sig <= to_unsigned(integer(my_rom(1963)),16);
when x"7ac" => lut_sig <= to_unsigned(integer(my_rom(1964)),16);
when x"7ad" => lut_sig <= to_unsigned(integer(my_rom(1965)),16);
when x"7ae" => lut_sig <= to_unsigned(integer(my_rom(1966)),16);
when x"7af" => lut_sig <= to_unsigned(integer(my_rom(1967)),16);
when x"7b0" => lut_sig <= to_unsigned(integer(my_rom(1968)),16);
when x"7b1" => lut_sig <= to_unsigned(integer(my_rom(1969)),16);
when x"7b2" => lut_sig <= to_unsigned(integer(my_rom(1970)),16);
when x"7b3" => lut_sig <= to_unsigned(integer(my_rom(1971)),16);
when x"7b4" => lut_sig <= to_unsigned(integer(my_rom(1972)),16);
when x"7b5" => lut_sig <= to_unsigned(integer(my_rom(1973)),16);
when x"7b6" => lut_sig <= to_unsigned(integer(my_rom(1974)),16);
when x"7b7" => lut_sig <= to_unsigned(integer(my_rom(1975)),16);
when x"7b8" => lut_sig <= to_unsigned(integer(my_rom(1976)),16);
when x"7b9" => lut_sig <= to_unsigned(integer(my_rom(1977)),16);
when x"7ba" => lut_sig <= to_unsigned(integer(my_rom(1978)),16);
when x"7bb" => lut_sig <= to_unsigned(integer(my_rom(1979)),16);
when x"7bc" => lut_sig <= to_unsigned(integer(my_rom(1980)),16);
when x"7bd" => lut_sig <= to_unsigned(integer(my_rom(1981)),16);
when x"7be" => lut_sig <= to_unsigned(integer(my_rom(1982)),16);
when x"7bf" => lut_sig <= to_unsigned(integer(my_rom(1983)),16);
when x"7c0" => lut_sig <= to_unsigned(integer(my_rom(1984)),16);
when x"7c1" => lut_sig <= to_unsigned(integer(my_rom(1985)),16);
when x"7c2" => lut_sig <= to_unsigned(integer(my_rom(1986)),16);
when x"7c3" => lut_sig <= to_unsigned(integer(my_rom(1987)),16);
when x"7c4" => lut_sig <= to_unsigned(integer(my_rom(1988)),16);
when x"7c5" => lut_sig <= to_unsigned(integer(my_rom(1989)),16);
when x"7c6" => lut_sig <= to_unsigned(integer(my_rom(1990)),16);
when x"7c7" => lut_sig <= to_unsigned(integer(my_rom(1991)),16);
when x"7c8" => lut_sig <= to_unsigned(integer(my_rom(1992)),16);
when x"7c9" => lut_sig <= to_unsigned(integer(my_rom(1993)),16);
when x"7ca" => lut_sig <= to_unsigned(integer(my_rom(1994)),16);
when x"7cb" => lut_sig <= to_unsigned(integer(my_rom(1995)),16);
when x"7cc" => lut_sig <= to_unsigned(integer(my_rom(1996)),16);
when x"7cd" => lut_sig <= to_unsigned(integer(my_rom(1997)),16);
when x"7ce" => lut_sig <= to_unsigned(integer(my_rom(1998)),16);
when x"7cf" => lut_sig <= to_unsigned(integer(my_rom(1999)),16);
when x"7d0" => lut_sig <= to_unsigned(integer(my_rom(2000)),16);
when x"7d1" => lut_sig <= to_unsigned(integer(my_rom(2001)),16);
when x"7d2" => lut_sig <= to_unsigned(integer(my_rom(2002)),16);
when x"7d3" => lut_sig <= to_unsigned(integer(my_rom(2003)),16);
when x"7d4" => lut_sig <= to_unsigned(integer(my_rom(2004)),16);
when x"7d5" => lut_sig <= to_unsigned(integer(my_rom(2005)),16);
when x"7d6" => lut_sig <= to_unsigned(integer(my_rom(2006)),16);
when x"7d7" => lut_sig <= to_unsigned(integer(my_rom(2007)),16);
when x"7d8" => lut_sig <= to_unsigned(integer(my_rom(2008)),16);
when x"7d9" => lut_sig <= to_unsigned(integer(my_rom(2009)),16);
when x"7da" => lut_sig <= to_unsigned(integer(my_rom(2010)),16);
when x"7db" => lut_sig <= to_unsigned(integer(my_rom(2011)),16);
when x"7dc" => lut_sig <= to_unsigned(integer(my_rom(2012)),16);
when x"7dd" => lut_sig <= to_unsigned(integer(my_rom(2013)),16);
when x"7de" => lut_sig <= to_unsigned(integer(my_rom(2014)),16);
when x"7df" => lut_sig <= to_unsigned(integer(my_rom(2015)),16);
when x"7e0" => lut_sig <= to_unsigned(integer(my_rom(2016)),16);
when x"7e1" => lut_sig <= to_unsigned(integer(my_rom(2017)),16);
when x"7e2" => lut_sig <= to_unsigned(integer(my_rom(2018)),16);
when x"7e3" => lut_sig <= to_unsigned(integer(my_rom(2019)),16);
when x"7e4" => lut_sig <= to_unsigned(integer(my_rom(2020)),16);
when x"7e5" => lut_sig <= to_unsigned(integer(my_rom(2021)),16);
when x"7e6" => lut_sig <= to_unsigned(integer(my_rom(2022)),16);
when x"7e7" => lut_sig <= to_unsigned(integer(my_rom(2023)),16);
when x"7e8" => lut_sig <= to_unsigned(integer(my_rom(2024)),16);
when x"7e9" => lut_sig <= to_unsigned(integer(my_rom(2025)),16);
when x"7ea" => lut_sig <= to_unsigned(integer(my_rom(2026)),16);
when x"7eb" => lut_sig <= to_unsigned(integer(my_rom(2027)),16);
when x"7ec" => lut_sig <= to_unsigned(integer(my_rom(2028)),16);
when x"7ed" => lut_sig <= to_unsigned(integer(my_rom(2029)),16);
when x"7ee" => lut_sig <= to_unsigned(integer(my_rom(2030)),16);
when x"7ef" => lut_sig <= to_unsigned(integer(my_rom(2031)),16);
when x"7f0" => lut_sig <= to_unsigned(integer(my_rom(2032)),16);
when x"7f1" => lut_sig <= to_unsigned(integer(my_rom(2033)),16);
when x"7f2" => lut_sig <= to_unsigned(integer(my_rom(2034)),16);
when x"7f3" => lut_sig <= to_unsigned(integer(my_rom(2035)),16);
when x"7f4" => lut_sig <= to_unsigned(integer(my_rom(2036)),16);
when x"7f5" => lut_sig <= to_unsigned(integer(my_rom(2037)),16);
when x"7f6" => lut_sig <= to_unsigned(integer(my_rom(2038)),16);
when x"7f7" => lut_sig <= to_unsigned(integer(my_rom(2039)),16);
when x"7f8" => lut_sig <= to_unsigned(integer(my_rom(2040)),16);
when x"7f9" => lut_sig <= to_unsigned(integer(my_rom(2041)),16);
when x"7fa" => lut_sig <= to_unsigned(integer(my_rom(2042)),16);
when x"7fb" => lut_sig <= to_unsigned(integer(my_rom(2043)),16);
when x"7fc" => lut_sig <= to_unsigned(integer(my_rom(2044)),16);
when x"7fd" => lut_sig <= to_unsigned(integer(my_rom(2045)),16);
when x"7fe" => lut_sig <= to_unsigned(integer(my_rom(2046)),16);
when x"7ff" => lut_sig <= to_unsigned(integer(my_rom(2047)),16);
when x"800" => lut_sig <= to_unsigned(integer(my_rom(2048)),16);
when x"801" => lut_sig <= to_unsigned(integer(my_rom(2049)),16);
when x"802" => lut_sig <= to_unsigned(integer(my_rom(2050)),16);
when x"803" => lut_sig <= to_unsigned(integer(my_rom(2051)),16);
when x"804" => lut_sig <= to_unsigned(integer(my_rom(2052)),16);
when x"805" => lut_sig <= to_unsigned(integer(my_rom(2053)),16);
when x"806" => lut_sig <= to_unsigned(integer(my_rom(2054)),16);
when x"807" => lut_sig <= to_unsigned(integer(my_rom(2055)),16);
when x"808" => lut_sig <= to_unsigned(integer(my_rom(2056)),16);
when x"809" => lut_sig <= to_unsigned(integer(my_rom(2057)),16);
when x"80a" => lut_sig <= to_unsigned(integer(my_rom(2058)),16);
when x"80b" => lut_sig <= to_unsigned(integer(my_rom(2059)),16);
when x"80c" => lut_sig <= to_unsigned(integer(my_rom(2060)),16);
when x"80d" => lut_sig <= to_unsigned(integer(my_rom(2061)),16);
when x"80e" => lut_sig <= to_unsigned(integer(my_rom(2062)),16);
when x"80f" => lut_sig <= to_unsigned(integer(my_rom(2063)),16);
when x"810" => lut_sig <= to_unsigned(integer(my_rom(2064)),16);
when x"811" => lut_sig <= to_unsigned(integer(my_rom(2065)),16);
when x"812" => lut_sig <= to_unsigned(integer(my_rom(2066)),16);
when x"813" => lut_sig <= to_unsigned(integer(my_rom(2067)),16);
when x"814" => lut_sig <= to_unsigned(integer(my_rom(2068)),16);
when x"815" => lut_sig <= to_unsigned(integer(my_rom(2069)),16);
when x"816" => lut_sig <= to_unsigned(integer(my_rom(2070)),16);
when x"817" => lut_sig <= to_unsigned(integer(my_rom(2071)),16);
when x"818" => lut_sig <= to_unsigned(integer(my_rom(2072)),16);
when x"819" => lut_sig <= to_unsigned(integer(my_rom(2073)),16);
when x"81a" => lut_sig <= to_unsigned(integer(my_rom(2074)),16);
when x"81b" => lut_sig <= to_unsigned(integer(my_rom(2075)),16);
when x"81c" => lut_sig <= to_unsigned(integer(my_rom(2076)),16);
when x"81d" => lut_sig <= to_unsigned(integer(my_rom(2077)),16);
when x"81e" => lut_sig <= to_unsigned(integer(my_rom(2078)),16);
when x"81f" => lut_sig <= to_unsigned(integer(my_rom(2079)),16);
when x"820" => lut_sig <= to_unsigned(integer(my_rom(2080)),16);
when x"821" => lut_sig <= to_unsigned(integer(my_rom(2081)),16);
when x"822" => lut_sig <= to_unsigned(integer(my_rom(2082)),16);
when x"823" => lut_sig <= to_unsigned(integer(my_rom(2083)),16);
when x"824" => lut_sig <= to_unsigned(integer(my_rom(2084)),16);
when x"825" => lut_sig <= to_unsigned(integer(my_rom(2085)),16);
when x"826" => lut_sig <= to_unsigned(integer(my_rom(2086)),16);
when x"827" => lut_sig <= to_unsigned(integer(my_rom(2087)),16);
when x"828" => lut_sig <= to_unsigned(integer(my_rom(2088)),16);
when x"829" => lut_sig <= to_unsigned(integer(my_rom(2089)),16);
when x"82a" => lut_sig <= to_unsigned(integer(my_rom(2090)),16);
when x"82b" => lut_sig <= to_unsigned(integer(my_rom(2091)),16);
when x"82c" => lut_sig <= to_unsigned(integer(my_rom(2092)),16);
when x"82d" => lut_sig <= to_unsigned(integer(my_rom(2093)),16);
when x"82e" => lut_sig <= to_unsigned(integer(my_rom(2094)),16);
when x"82f" => lut_sig <= to_unsigned(integer(my_rom(2095)),16);
when x"830" => lut_sig <= to_unsigned(integer(my_rom(2096)),16);
when x"831" => lut_sig <= to_unsigned(integer(my_rom(2097)),16);
when x"832" => lut_sig <= to_unsigned(integer(my_rom(2098)),16);
when x"833" => lut_sig <= to_unsigned(integer(my_rom(2099)),16);
when x"834" => lut_sig <= to_unsigned(integer(my_rom(2100)),16);
when x"835" => lut_sig <= to_unsigned(integer(my_rom(2101)),16);
when x"836" => lut_sig <= to_unsigned(integer(my_rom(2102)),16);
when x"837" => lut_sig <= to_unsigned(integer(my_rom(2103)),16);
when x"838" => lut_sig <= to_unsigned(integer(my_rom(2104)),16);
when x"839" => lut_sig <= to_unsigned(integer(my_rom(2105)),16);
when x"83a" => lut_sig <= to_unsigned(integer(my_rom(2106)),16);
when x"83b" => lut_sig <= to_unsigned(integer(my_rom(2107)),16);
when x"83c" => lut_sig <= to_unsigned(integer(my_rom(2108)),16);
when x"83d" => lut_sig <= to_unsigned(integer(my_rom(2109)),16);
when x"83e" => lut_sig <= to_unsigned(integer(my_rom(2110)),16);
when x"83f" => lut_sig <= to_unsigned(integer(my_rom(2111)),16);
when x"840" => lut_sig <= to_unsigned(integer(my_rom(2112)),16);
when x"841" => lut_sig <= to_unsigned(integer(my_rom(2113)),16);
when x"842" => lut_sig <= to_unsigned(integer(my_rom(2114)),16);
when x"843" => lut_sig <= to_unsigned(integer(my_rom(2115)),16);
when x"844" => lut_sig <= to_unsigned(integer(my_rom(2116)),16);
when x"845" => lut_sig <= to_unsigned(integer(my_rom(2117)),16);
when x"846" => lut_sig <= to_unsigned(integer(my_rom(2118)),16);
when x"847" => lut_sig <= to_unsigned(integer(my_rom(2119)),16);
when x"848" => lut_sig <= to_unsigned(integer(my_rom(2120)),16);
when x"849" => lut_sig <= to_unsigned(integer(my_rom(2121)),16);
when x"84a" => lut_sig <= to_unsigned(integer(my_rom(2122)),16);
when x"84b" => lut_sig <= to_unsigned(integer(my_rom(2123)),16);
when x"84c" => lut_sig <= to_unsigned(integer(my_rom(2124)),16);
when x"84d" => lut_sig <= to_unsigned(integer(my_rom(2125)),16);
when x"84e" => lut_sig <= to_unsigned(integer(my_rom(2126)),16);
when x"84f" => lut_sig <= to_unsigned(integer(my_rom(2127)),16);
when x"850" => lut_sig <= to_unsigned(integer(my_rom(2128)),16);
when x"851" => lut_sig <= to_unsigned(integer(my_rom(2129)),16);
when x"852" => lut_sig <= to_unsigned(integer(my_rom(2130)),16);
when x"853" => lut_sig <= to_unsigned(integer(my_rom(2131)),16);
when x"854" => lut_sig <= to_unsigned(integer(my_rom(2132)),16);
when x"855" => lut_sig <= to_unsigned(integer(my_rom(2133)),16);
when x"856" => lut_sig <= to_unsigned(integer(my_rom(2134)),16);
when x"857" => lut_sig <= to_unsigned(integer(my_rom(2135)),16);
when x"858" => lut_sig <= to_unsigned(integer(my_rom(2136)),16);
when x"859" => lut_sig <= to_unsigned(integer(my_rom(2137)),16);
when x"85a" => lut_sig <= to_unsigned(integer(my_rom(2138)),16);
when x"85b" => lut_sig <= to_unsigned(integer(my_rom(2139)),16);
when x"85c" => lut_sig <= to_unsigned(integer(my_rom(2140)),16);
when x"85d" => lut_sig <= to_unsigned(integer(my_rom(2141)),16);
when x"85e" => lut_sig <= to_unsigned(integer(my_rom(2142)),16);
when x"85f" => lut_sig <= to_unsigned(integer(my_rom(2143)),16);
when x"860" => lut_sig <= to_unsigned(integer(my_rom(2144)),16);
when x"861" => lut_sig <= to_unsigned(integer(my_rom(2145)),16);
when x"862" => lut_sig <= to_unsigned(integer(my_rom(2146)),16);
when x"863" => lut_sig <= to_unsigned(integer(my_rom(2147)),16);
when x"864" => lut_sig <= to_unsigned(integer(my_rom(2148)),16);
when x"865" => lut_sig <= to_unsigned(integer(my_rom(2149)),16);
when x"866" => lut_sig <= to_unsigned(integer(my_rom(2150)),16);
when x"867" => lut_sig <= to_unsigned(integer(my_rom(2151)),16);
when x"868" => lut_sig <= to_unsigned(integer(my_rom(2152)),16);
when x"869" => lut_sig <= to_unsigned(integer(my_rom(2153)),16);
when x"86a" => lut_sig <= to_unsigned(integer(my_rom(2154)),16);
when x"86b" => lut_sig <= to_unsigned(integer(my_rom(2155)),16);
when x"86c" => lut_sig <= to_unsigned(integer(my_rom(2156)),16);
when x"86d" => lut_sig <= to_unsigned(integer(my_rom(2157)),16);
when x"86e" => lut_sig <= to_unsigned(integer(my_rom(2158)),16);
when x"86f" => lut_sig <= to_unsigned(integer(my_rom(2159)),16);
when x"870" => lut_sig <= to_unsigned(integer(my_rom(2160)),16);
when x"871" => lut_sig <= to_unsigned(integer(my_rom(2161)),16);
when x"872" => lut_sig <= to_unsigned(integer(my_rom(2162)),16);
when x"873" => lut_sig <= to_unsigned(integer(my_rom(2163)),16);
when x"874" => lut_sig <= to_unsigned(integer(my_rom(2164)),16);
when x"875" => lut_sig <= to_unsigned(integer(my_rom(2165)),16);
when x"876" => lut_sig <= to_unsigned(integer(my_rom(2166)),16);
when x"877" => lut_sig <= to_unsigned(integer(my_rom(2167)),16);
when x"878" => lut_sig <= to_unsigned(integer(my_rom(2168)),16);
when x"879" => lut_sig <= to_unsigned(integer(my_rom(2169)),16);
when x"87a" => lut_sig <= to_unsigned(integer(my_rom(2170)),16);
when x"87b" => lut_sig <= to_unsigned(integer(my_rom(2171)),16);
when x"87c" => lut_sig <= to_unsigned(integer(my_rom(2172)),16);
when x"87d" => lut_sig <= to_unsigned(integer(my_rom(2173)),16);
when x"87e" => lut_sig <= to_unsigned(integer(my_rom(2174)),16);
when x"87f" => lut_sig <= to_unsigned(integer(my_rom(2175)),16);
when x"880" => lut_sig <= to_unsigned(integer(my_rom(2176)),16);
when x"881" => lut_sig <= to_unsigned(integer(my_rom(2177)),16);
when x"882" => lut_sig <= to_unsigned(integer(my_rom(2178)),16);
when x"883" => lut_sig <= to_unsigned(integer(my_rom(2179)),16);
when x"884" => lut_sig <= to_unsigned(integer(my_rom(2180)),16);
when x"885" => lut_sig <= to_unsigned(integer(my_rom(2181)),16);
when x"886" => lut_sig <= to_unsigned(integer(my_rom(2182)),16);
when x"887" => lut_sig <= to_unsigned(integer(my_rom(2183)),16);
when x"888" => lut_sig <= to_unsigned(integer(my_rom(2184)),16);
when x"889" => lut_sig <= to_unsigned(integer(my_rom(2185)),16);
when x"88a" => lut_sig <= to_unsigned(integer(my_rom(2186)),16);
when x"88b" => lut_sig <= to_unsigned(integer(my_rom(2187)),16);
when x"88c" => lut_sig <= to_unsigned(integer(my_rom(2188)),16);
when x"88d" => lut_sig <= to_unsigned(integer(my_rom(2189)),16);
when x"88e" => lut_sig <= to_unsigned(integer(my_rom(2190)),16);
when x"88f" => lut_sig <= to_unsigned(integer(my_rom(2191)),16);
when x"890" => lut_sig <= to_unsigned(integer(my_rom(2192)),16);
when x"891" => lut_sig <= to_unsigned(integer(my_rom(2193)),16);
when x"892" => lut_sig <= to_unsigned(integer(my_rom(2194)),16);
when x"893" => lut_sig <= to_unsigned(integer(my_rom(2195)),16);
when x"894" => lut_sig <= to_unsigned(integer(my_rom(2196)),16);
when x"895" => lut_sig <= to_unsigned(integer(my_rom(2197)),16);
when x"896" => lut_sig <= to_unsigned(integer(my_rom(2198)),16);
when x"897" => lut_sig <= to_unsigned(integer(my_rom(2199)),16);
when x"898" => lut_sig <= to_unsigned(integer(my_rom(2200)),16);
when x"899" => lut_sig <= to_unsigned(integer(my_rom(2201)),16);
when x"89a" => lut_sig <= to_unsigned(integer(my_rom(2202)),16);
when x"89b" => lut_sig <= to_unsigned(integer(my_rom(2203)),16);
when x"89c" => lut_sig <= to_unsigned(integer(my_rom(2204)),16);
when x"89d" => lut_sig <= to_unsigned(integer(my_rom(2205)),16);
when x"89e" => lut_sig <= to_unsigned(integer(my_rom(2206)),16);
when x"89f" => lut_sig <= to_unsigned(integer(my_rom(2207)),16);
when x"8a0" => lut_sig <= to_unsigned(integer(my_rom(2208)),16);
when x"8a1" => lut_sig <= to_unsigned(integer(my_rom(2209)),16);
when x"8a2" => lut_sig <= to_unsigned(integer(my_rom(2210)),16);
when x"8a3" => lut_sig <= to_unsigned(integer(my_rom(2211)),16);
when x"8a4" => lut_sig <= to_unsigned(integer(my_rom(2212)),16);
when x"8a5" => lut_sig <= to_unsigned(integer(my_rom(2213)),16);
when x"8a6" => lut_sig <= to_unsigned(integer(my_rom(2214)),16);
when x"8a7" => lut_sig <= to_unsigned(integer(my_rom(2215)),16);
when x"8a8" => lut_sig <= to_unsigned(integer(my_rom(2216)),16);
when x"8a9" => lut_sig <= to_unsigned(integer(my_rom(2217)),16);
when x"8aa" => lut_sig <= to_unsigned(integer(my_rom(2218)),16);
when x"8ab" => lut_sig <= to_unsigned(integer(my_rom(2219)),16);
when x"8ac" => lut_sig <= to_unsigned(integer(my_rom(2220)),16);
when x"8ad" => lut_sig <= to_unsigned(integer(my_rom(2221)),16);
when x"8ae" => lut_sig <= to_unsigned(integer(my_rom(2222)),16);
when x"8af" => lut_sig <= to_unsigned(integer(my_rom(2223)),16);
when x"8b0" => lut_sig <= to_unsigned(integer(my_rom(2224)),16);
when x"8b1" => lut_sig <= to_unsigned(integer(my_rom(2225)),16);
when x"8b2" => lut_sig <= to_unsigned(integer(my_rom(2226)),16);
when x"8b3" => lut_sig <= to_unsigned(integer(my_rom(2227)),16);
when x"8b4" => lut_sig <= to_unsigned(integer(my_rom(2228)),16);
when x"8b5" => lut_sig <= to_unsigned(integer(my_rom(2229)),16);
when x"8b6" => lut_sig <= to_unsigned(integer(my_rom(2230)),16);
when x"8b7" => lut_sig <= to_unsigned(integer(my_rom(2231)),16);
when x"8b8" => lut_sig <= to_unsigned(integer(my_rom(2232)),16);
when x"8b9" => lut_sig <= to_unsigned(integer(my_rom(2233)),16);
when x"8ba" => lut_sig <= to_unsigned(integer(my_rom(2234)),16);
when x"8bb" => lut_sig <= to_unsigned(integer(my_rom(2235)),16);
when x"8bc" => lut_sig <= to_unsigned(integer(my_rom(2236)),16);
when x"8bd" => lut_sig <= to_unsigned(integer(my_rom(2237)),16);
when x"8be" => lut_sig <= to_unsigned(integer(my_rom(2238)),16);
when x"8bf" => lut_sig <= to_unsigned(integer(my_rom(2239)),16);
when x"8c0" => lut_sig <= to_unsigned(integer(my_rom(2240)),16);
when x"8c1" => lut_sig <= to_unsigned(integer(my_rom(2241)),16);
when x"8c2" => lut_sig <= to_unsigned(integer(my_rom(2242)),16);
when x"8c3" => lut_sig <= to_unsigned(integer(my_rom(2243)),16);
when x"8c4" => lut_sig <= to_unsigned(integer(my_rom(2244)),16);
when x"8c5" => lut_sig <= to_unsigned(integer(my_rom(2245)),16);
when x"8c6" => lut_sig <= to_unsigned(integer(my_rom(2246)),16);
when x"8c7" => lut_sig <= to_unsigned(integer(my_rom(2247)),16);
when x"8c8" => lut_sig <= to_unsigned(integer(my_rom(2248)),16);
when x"8c9" => lut_sig <= to_unsigned(integer(my_rom(2249)),16);
when x"8ca" => lut_sig <= to_unsigned(integer(my_rom(2250)),16);
when x"8cb" => lut_sig <= to_unsigned(integer(my_rom(2251)),16);
when x"8cc" => lut_sig <= to_unsigned(integer(my_rom(2252)),16);
when x"8cd" => lut_sig <= to_unsigned(integer(my_rom(2253)),16);
when x"8ce" => lut_sig <= to_unsigned(integer(my_rom(2254)),16);
when x"8cf" => lut_sig <= to_unsigned(integer(my_rom(2255)),16);
when x"8d0" => lut_sig <= to_unsigned(integer(my_rom(2256)),16);
when x"8d1" => lut_sig <= to_unsigned(integer(my_rom(2257)),16);
when x"8d2" => lut_sig <= to_unsigned(integer(my_rom(2258)),16);
when x"8d3" => lut_sig <= to_unsigned(integer(my_rom(2259)),16);
when x"8d4" => lut_sig <= to_unsigned(integer(my_rom(2260)),16);
when x"8d5" => lut_sig <= to_unsigned(integer(my_rom(2261)),16);
when x"8d6" => lut_sig <= to_unsigned(integer(my_rom(2262)),16);
when x"8d7" => lut_sig <= to_unsigned(integer(my_rom(2263)),16);
when x"8d8" => lut_sig <= to_unsigned(integer(my_rom(2264)),16);
when x"8d9" => lut_sig <= to_unsigned(integer(my_rom(2265)),16);
when x"8da" => lut_sig <= to_unsigned(integer(my_rom(2266)),16);
when x"8db" => lut_sig <= to_unsigned(integer(my_rom(2267)),16);
when x"8dc" => lut_sig <= to_unsigned(integer(my_rom(2268)),16);
when x"8dd" => lut_sig <= to_unsigned(integer(my_rom(2269)),16);
when x"8de" => lut_sig <= to_unsigned(integer(my_rom(2270)),16);
when x"8df" => lut_sig <= to_unsigned(integer(my_rom(2271)),16);
when x"8e0" => lut_sig <= to_unsigned(integer(my_rom(2272)),16);
when x"8e1" => lut_sig <= to_unsigned(integer(my_rom(2273)),16);
when x"8e2" => lut_sig <= to_unsigned(integer(my_rom(2274)),16);
when x"8e3" => lut_sig <= to_unsigned(integer(my_rom(2275)),16);
when x"8e4" => lut_sig <= to_unsigned(integer(my_rom(2276)),16);
when x"8e5" => lut_sig <= to_unsigned(integer(my_rom(2277)),16);
when x"8e6" => lut_sig <= to_unsigned(integer(my_rom(2278)),16);
when x"8e7" => lut_sig <= to_unsigned(integer(my_rom(2279)),16);
when x"8e8" => lut_sig <= to_unsigned(integer(my_rom(2280)),16);
when x"8e9" => lut_sig <= to_unsigned(integer(my_rom(2281)),16);
when x"8ea" => lut_sig <= to_unsigned(integer(my_rom(2282)),16);
when x"8eb" => lut_sig <= to_unsigned(integer(my_rom(2283)),16);
when x"8ec" => lut_sig <= to_unsigned(integer(my_rom(2284)),16);
when x"8ed" => lut_sig <= to_unsigned(integer(my_rom(2285)),16);
when x"8ee" => lut_sig <= to_unsigned(integer(my_rom(2286)),16);
when x"8ef" => lut_sig <= to_unsigned(integer(my_rom(2287)),16);
when x"8f0" => lut_sig <= to_unsigned(integer(my_rom(2288)),16);
when x"8f1" => lut_sig <= to_unsigned(integer(my_rom(2289)),16);
when x"8f2" => lut_sig <= to_unsigned(integer(my_rom(2290)),16);
when x"8f3" => lut_sig <= to_unsigned(integer(my_rom(2291)),16);
when x"8f4" => lut_sig <= to_unsigned(integer(my_rom(2292)),16);
when x"8f5" => lut_sig <= to_unsigned(integer(my_rom(2293)),16);
when x"8f6" => lut_sig <= to_unsigned(integer(my_rom(2294)),16);
when x"8f7" => lut_sig <= to_unsigned(integer(my_rom(2295)),16);
when x"8f8" => lut_sig <= to_unsigned(integer(my_rom(2296)),16);
when x"8f9" => lut_sig <= to_unsigned(integer(my_rom(2297)),16);
when x"8fa" => lut_sig <= to_unsigned(integer(my_rom(2298)),16);
when x"8fb" => lut_sig <= to_unsigned(integer(my_rom(2299)),16);
when x"8fc" => lut_sig <= to_unsigned(integer(my_rom(2300)),16);
when x"8fd" => lut_sig <= to_unsigned(integer(my_rom(2301)),16);
when x"8fe" => lut_sig <= to_unsigned(integer(my_rom(2302)),16);
when x"8ff" => lut_sig <= to_unsigned(integer(my_rom(2303)),16);
when x"900" => lut_sig <= to_unsigned(integer(my_rom(2304)),16);
when x"901" => lut_sig <= to_unsigned(integer(my_rom(2305)),16);
when x"902" => lut_sig <= to_unsigned(integer(my_rom(2306)),16);
when x"903" => lut_sig <= to_unsigned(integer(my_rom(2307)),16);
when x"904" => lut_sig <= to_unsigned(integer(my_rom(2308)),16);
when x"905" => lut_sig <= to_unsigned(integer(my_rom(2309)),16);
when x"906" => lut_sig <= to_unsigned(integer(my_rom(2310)),16);
when x"907" => lut_sig <= to_unsigned(integer(my_rom(2311)),16);
when x"908" => lut_sig <= to_unsigned(integer(my_rom(2312)),16);
when x"909" => lut_sig <= to_unsigned(integer(my_rom(2313)),16);
when x"90a" => lut_sig <= to_unsigned(integer(my_rom(2314)),16);
when x"90b" => lut_sig <= to_unsigned(integer(my_rom(2315)),16);
when x"90c" => lut_sig <= to_unsigned(integer(my_rom(2316)),16);
when x"90d" => lut_sig <= to_unsigned(integer(my_rom(2317)),16);
when x"90e" => lut_sig <= to_unsigned(integer(my_rom(2318)),16);
when x"90f" => lut_sig <= to_unsigned(integer(my_rom(2319)),16);
when x"910" => lut_sig <= to_unsigned(integer(my_rom(2320)),16);
when x"911" => lut_sig <= to_unsigned(integer(my_rom(2321)),16);
when x"912" => lut_sig <= to_unsigned(integer(my_rom(2322)),16);
when x"913" => lut_sig <= to_unsigned(integer(my_rom(2323)),16);
when x"914" => lut_sig <= to_unsigned(integer(my_rom(2324)),16);
when x"915" => lut_sig <= to_unsigned(integer(my_rom(2325)),16);
when x"916" => lut_sig <= to_unsigned(integer(my_rom(2326)),16);
when x"917" => lut_sig <= to_unsigned(integer(my_rom(2327)),16);
when x"918" => lut_sig <= to_unsigned(integer(my_rom(2328)),16);
when x"919" => lut_sig <= to_unsigned(integer(my_rom(2329)),16);
when x"91a" => lut_sig <= to_unsigned(integer(my_rom(2330)),16);
when x"91b" => lut_sig <= to_unsigned(integer(my_rom(2331)),16);
when x"91c" => lut_sig <= to_unsigned(integer(my_rom(2332)),16);
when x"91d" => lut_sig <= to_unsigned(integer(my_rom(2333)),16);
when x"91e" => lut_sig <= to_unsigned(integer(my_rom(2334)),16);
when x"91f" => lut_sig <= to_unsigned(integer(my_rom(2335)),16);
when x"920" => lut_sig <= to_unsigned(integer(my_rom(2336)),16);
when x"921" => lut_sig <= to_unsigned(integer(my_rom(2337)),16);
when x"922" => lut_sig <= to_unsigned(integer(my_rom(2338)),16);
when x"923" => lut_sig <= to_unsigned(integer(my_rom(2339)),16);
when x"924" => lut_sig <= to_unsigned(integer(my_rom(2340)),16);
when x"925" => lut_sig <= to_unsigned(integer(my_rom(2341)),16);
when x"926" => lut_sig <= to_unsigned(integer(my_rom(2342)),16);
when x"927" => lut_sig <= to_unsigned(integer(my_rom(2343)),16);
when x"928" => lut_sig <= to_unsigned(integer(my_rom(2344)),16);
when x"929" => lut_sig <= to_unsigned(integer(my_rom(2345)),16);
when x"92a" => lut_sig <= to_unsigned(integer(my_rom(2346)),16);
when x"92b" => lut_sig <= to_unsigned(integer(my_rom(2347)),16);
when x"92c" => lut_sig <= to_unsigned(integer(my_rom(2348)),16);
when x"92d" => lut_sig <= to_unsigned(integer(my_rom(2349)),16);
when x"92e" => lut_sig <= to_unsigned(integer(my_rom(2350)),16);
when x"92f" => lut_sig <= to_unsigned(integer(my_rom(2351)),16);
when x"930" => lut_sig <= to_unsigned(integer(my_rom(2352)),16);
when x"931" => lut_sig <= to_unsigned(integer(my_rom(2353)),16);
when x"932" => lut_sig <= to_unsigned(integer(my_rom(2354)),16);
when x"933" => lut_sig <= to_unsigned(integer(my_rom(2355)),16);
when x"934" => lut_sig <= to_unsigned(integer(my_rom(2356)),16);
when x"935" => lut_sig <= to_unsigned(integer(my_rom(2357)),16);
when x"936" => lut_sig <= to_unsigned(integer(my_rom(2358)),16);
when x"937" => lut_sig <= to_unsigned(integer(my_rom(2359)),16);
when x"938" => lut_sig <= to_unsigned(integer(my_rom(2360)),16);
when x"939" => lut_sig <= to_unsigned(integer(my_rom(2361)),16);
when x"93a" => lut_sig <= to_unsigned(integer(my_rom(2362)),16);
when x"93b" => lut_sig <= to_unsigned(integer(my_rom(2363)),16);
when x"93c" => lut_sig <= to_unsigned(integer(my_rom(2364)),16);
when x"93d" => lut_sig <= to_unsigned(integer(my_rom(2365)),16);
when x"93e" => lut_sig <= to_unsigned(integer(my_rom(2366)),16);
when x"93f" => lut_sig <= to_unsigned(integer(my_rom(2367)),16);
when x"940" => lut_sig <= to_unsigned(integer(my_rom(2368)),16);
when x"941" => lut_sig <= to_unsigned(integer(my_rom(2369)),16);
when x"942" => lut_sig <= to_unsigned(integer(my_rom(2370)),16);
when x"943" => lut_sig <= to_unsigned(integer(my_rom(2371)),16);
when x"944" => lut_sig <= to_unsigned(integer(my_rom(2372)),16);
when x"945" => lut_sig <= to_unsigned(integer(my_rom(2373)),16);
when x"946" => lut_sig <= to_unsigned(integer(my_rom(2374)),16);
when x"947" => lut_sig <= to_unsigned(integer(my_rom(2375)),16);
when x"948" => lut_sig <= to_unsigned(integer(my_rom(2376)),16);
when x"949" => lut_sig <= to_unsigned(integer(my_rom(2377)),16);
when x"94a" => lut_sig <= to_unsigned(integer(my_rom(2378)),16);
when x"94b" => lut_sig <= to_unsigned(integer(my_rom(2379)),16);
when x"94c" => lut_sig <= to_unsigned(integer(my_rom(2380)),16);
when x"94d" => lut_sig <= to_unsigned(integer(my_rom(2381)),16);
when x"94e" => lut_sig <= to_unsigned(integer(my_rom(2382)),16);
when x"94f" => lut_sig <= to_unsigned(integer(my_rom(2383)),16);
when x"950" => lut_sig <= to_unsigned(integer(my_rom(2384)),16);
when x"951" => lut_sig <= to_unsigned(integer(my_rom(2385)),16);
when x"952" => lut_sig <= to_unsigned(integer(my_rom(2386)),16);
when x"953" => lut_sig <= to_unsigned(integer(my_rom(2387)),16);
when x"954" => lut_sig <= to_unsigned(integer(my_rom(2388)),16);
when x"955" => lut_sig <= to_unsigned(integer(my_rom(2389)),16);
when x"956" => lut_sig <= to_unsigned(integer(my_rom(2390)),16);
when x"957" => lut_sig <= to_unsigned(integer(my_rom(2391)),16);
when x"958" => lut_sig <= to_unsigned(integer(my_rom(2392)),16);
when x"959" => lut_sig <= to_unsigned(integer(my_rom(2393)),16);
when x"95a" => lut_sig <= to_unsigned(integer(my_rom(2394)),16);
when x"95b" => lut_sig <= to_unsigned(integer(my_rom(2395)),16);
when x"95c" => lut_sig <= to_unsigned(integer(my_rom(2396)),16);
when x"95d" => lut_sig <= to_unsigned(integer(my_rom(2397)),16);
when x"95e" => lut_sig <= to_unsigned(integer(my_rom(2398)),16);
when x"95f" => lut_sig <= to_unsigned(integer(my_rom(2399)),16);
when x"960" => lut_sig <= to_unsigned(integer(my_rom(2400)),16);
when x"961" => lut_sig <= to_unsigned(integer(my_rom(2401)),16);
when x"962" => lut_sig <= to_unsigned(integer(my_rom(2402)),16);
when x"963" => lut_sig <= to_unsigned(integer(my_rom(2403)),16);
when x"964" => lut_sig <= to_unsigned(integer(my_rom(2404)),16);
when x"965" => lut_sig <= to_unsigned(integer(my_rom(2405)),16);
when x"966" => lut_sig <= to_unsigned(integer(my_rom(2406)),16);
when x"967" => lut_sig <= to_unsigned(integer(my_rom(2407)),16);
when x"968" => lut_sig <= to_unsigned(integer(my_rom(2408)),16);
when x"969" => lut_sig <= to_unsigned(integer(my_rom(2409)),16);
when x"96a" => lut_sig <= to_unsigned(integer(my_rom(2410)),16);
when x"96b" => lut_sig <= to_unsigned(integer(my_rom(2411)),16);
when x"96c" => lut_sig <= to_unsigned(integer(my_rom(2412)),16);
when x"96d" => lut_sig <= to_unsigned(integer(my_rom(2413)),16);
when x"96e" => lut_sig <= to_unsigned(integer(my_rom(2414)),16);
when x"96f" => lut_sig <= to_unsigned(integer(my_rom(2415)),16);
when x"970" => lut_sig <= to_unsigned(integer(my_rom(2416)),16);
when x"971" => lut_sig <= to_unsigned(integer(my_rom(2417)),16);
when x"972" => lut_sig <= to_unsigned(integer(my_rom(2418)),16);
when x"973" => lut_sig <= to_unsigned(integer(my_rom(2419)),16);
when x"974" => lut_sig <= to_unsigned(integer(my_rom(2420)),16);
when x"975" => lut_sig <= to_unsigned(integer(my_rom(2421)),16);
when x"976" => lut_sig <= to_unsigned(integer(my_rom(2422)),16);
when x"977" => lut_sig <= to_unsigned(integer(my_rom(2423)),16);
when x"978" => lut_sig <= to_unsigned(integer(my_rom(2424)),16);
when x"979" => lut_sig <= to_unsigned(integer(my_rom(2425)),16);
when x"97a" => lut_sig <= to_unsigned(integer(my_rom(2426)),16);
when x"97b" => lut_sig <= to_unsigned(integer(my_rom(2427)),16);
when x"97c" => lut_sig <= to_unsigned(integer(my_rom(2428)),16);
when x"97d" => lut_sig <= to_unsigned(integer(my_rom(2429)),16);
when x"97e" => lut_sig <= to_unsigned(integer(my_rom(2430)),16);
when x"97f" => lut_sig <= to_unsigned(integer(my_rom(2431)),16);
when x"980" => lut_sig <= to_unsigned(integer(my_rom(2432)),16);
when x"981" => lut_sig <= to_unsigned(integer(my_rom(2433)),16);
when x"982" => lut_sig <= to_unsigned(integer(my_rom(2434)),16);
when x"983" => lut_sig <= to_unsigned(integer(my_rom(2435)),16);
when x"984" => lut_sig <= to_unsigned(integer(my_rom(2436)),16);
when x"985" => lut_sig <= to_unsigned(integer(my_rom(2437)),16);
when x"986" => lut_sig <= to_unsigned(integer(my_rom(2438)),16);
when x"987" => lut_sig <= to_unsigned(integer(my_rom(2439)),16);
when x"988" => lut_sig <= to_unsigned(integer(my_rom(2440)),16);
when x"989" => lut_sig <= to_unsigned(integer(my_rom(2441)),16);
when x"98a" => lut_sig <= to_unsigned(integer(my_rom(2442)),16);
when x"98b" => lut_sig <= to_unsigned(integer(my_rom(2443)),16);
when x"98c" => lut_sig <= to_unsigned(integer(my_rom(2444)),16);
when x"98d" => lut_sig <= to_unsigned(integer(my_rom(2445)),16);
when x"98e" => lut_sig <= to_unsigned(integer(my_rom(2446)),16);
when x"98f" => lut_sig <= to_unsigned(integer(my_rom(2447)),16);
when x"990" => lut_sig <= to_unsigned(integer(my_rom(2448)),16);
when x"991" => lut_sig <= to_unsigned(integer(my_rom(2449)),16);
when x"992" => lut_sig <= to_unsigned(integer(my_rom(2450)),16);
when x"993" => lut_sig <= to_unsigned(integer(my_rom(2451)),16);
when x"994" => lut_sig <= to_unsigned(integer(my_rom(2452)),16);
when x"995" => lut_sig <= to_unsigned(integer(my_rom(2453)),16);
when x"996" => lut_sig <= to_unsigned(integer(my_rom(2454)),16);
when x"997" => lut_sig <= to_unsigned(integer(my_rom(2455)),16);
when x"998" => lut_sig <= to_unsigned(integer(my_rom(2456)),16);
when x"999" => lut_sig <= to_unsigned(integer(my_rom(2457)),16);
when x"99a" => lut_sig <= to_unsigned(integer(my_rom(2458)),16);
when x"99b" => lut_sig <= to_unsigned(integer(my_rom(2459)),16);
when x"99c" => lut_sig <= to_unsigned(integer(my_rom(2460)),16);
when x"99d" => lut_sig <= to_unsigned(integer(my_rom(2461)),16);
when x"99e" => lut_sig <= to_unsigned(integer(my_rom(2462)),16);
when x"99f" => lut_sig <= to_unsigned(integer(my_rom(2463)),16);
when x"9a0" => lut_sig <= to_unsigned(integer(my_rom(2464)),16);
when x"9a1" => lut_sig <= to_unsigned(integer(my_rom(2465)),16);
when x"9a2" => lut_sig <= to_unsigned(integer(my_rom(2466)),16);
when x"9a3" => lut_sig <= to_unsigned(integer(my_rom(2467)),16);
when x"9a4" => lut_sig <= to_unsigned(integer(my_rom(2468)),16);
when x"9a5" => lut_sig <= to_unsigned(integer(my_rom(2469)),16);
when x"9a6" => lut_sig <= to_unsigned(integer(my_rom(2470)),16);
when x"9a7" => lut_sig <= to_unsigned(integer(my_rom(2471)),16);
when x"9a8" => lut_sig <= to_unsigned(integer(my_rom(2472)),16);
when x"9a9" => lut_sig <= to_unsigned(integer(my_rom(2473)),16);
when x"9aa" => lut_sig <= to_unsigned(integer(my_rom(2474)),16);
when x"9ab" => lut_sig <= to_unsigned(integer(my_rom(2475)),16);
when x"9ac" => lut_sig <= to_unsigned(integer(my_rom(2476)),16);
when x"9ad" => lut_sig <= to_unsigned(integer(my_rom(2477)),16);
when x"9ae" => lut_sig <= to_unsigned(integer(my_rom(2478)),16);
when x"9af" => lut_sig <= to_unsigned(integer(my_rom(2479)),16);
when x"9b0" => lut_sig <= to_unsigned(integer(my_rom(2480)),16);
when x"9b1" => lut_sig <= to_unsigned(integer(my_rom(2481)),16);
when x"9b2" => lut_sig <= to_unsigned(integer(my_rom(2482)),16);
when x"9b3" => lut_sig <= to_unsigned(integer(my_rom(2483)),16);
when x"9b4" => lut_sig <= to_unsigned(integer(my_rom(2484)),16);
when x"9b5" => lut_sig <= to_unsigned(integer(my_rom(2485)),16);
when x"9b6" => lut_sig <= to_unsigned(integer(my_rom(2486)),16);
when x"9b7" => lut_sig <= to_unsigned(integer(my_rom(2487)),16);
when x"9b8" => lut_sig <= to_unsigned(integer(my_rom(2488)),16);
when x"9b9" => lut_sig <= to_unsigned(integer(my_rom(2489)),16);
when x"9ba" => lut_sig <= to_unsigned(integer(my_rom(2490)),16);
when x"9bb" => lut_sig <= to_unsigned(integer(my_rom(2491)),16);
when x"9bc" => lut_sig <= to_unsigned(integer(my_rom(2492)),16);
when x"9bd" => lut_sig <= to_unsigned(integer(my_rom(2493)),16);
when x"9be" => lut_sig <= to_unsigned(integer(my_rom(2494)),16);
when x"9bf" => lut_sig <= to_unsigned(integer(my_rom(2495)),16);
when x"9c0" => lut_sig <= to_unsigned(integer(my_rom(2496)),16);
when x"9c1" => lut_sig <= to_unsigned(integer(my_rom(2497)),16);
when x"9c2" => lut_sig <= to_unsigned(integer(my_rom(2498)),16);
when x"9c3" => lut_sig <= to_unsigned(integer(my_rom(2499)),16);
when x"9c4" => lut_sig <= to_unsigned(integer(my_rom(2500)),16);
when x"9c5" => lut_sig <= to_unsigned(integer(my_rom(2501)),16);
when x"9c6" => lut_sig <= to_unsigned(integer(my_rom(2502)),16);
when x"9c7" => lut_sig <= to_unsigned(integer(my_rom(2503)),16);
when x"9c8" => lut_sig <= to_unsigned(integer(my_rom(2504)),16);
when x"9c9" => lut_sig <= to_unsigned(integer(my_rom(2505)),16);
when x"9ca" => lut_sig <= to_unsigned(integer(my_rom(2506)),16);
when x"9cb" => lut_sig <= to_unsigned(integer(my_rom(2507)),16);
when x"9cc" => lut_sig <= to_unsigned(integer(my_rom(2508)),16);
when x"9cd" => lut_sig <= to_unsigned(integer(my_rom(2509)),16);
when x"9ce" => lut_sig <= to_unsigned(integer(my_rom(2510)),16);
when x"9cf" => lut_sig <= to_unsigned(integer(my_rom(2511)),16);
when x"9d0" => lut_sig <= to_unsigned(integer(my_rom(2512)),16);
when x"9d1" => lut_sig <= to_unsigned(integer(my_rom(2513)),16);
when x"9d2" => lut_sig <= to_unsigned(integer(my_rom(2514)),16);
when x"9d3" => lut_sig <= to_unsigned(integer(my_rom(2515)),16);
when x"9d4" => lut_sig <= to_unsigned(integer(my_rom(2516)),16);
when x"9d5" => lut_sig <= to_unsigned(integer(my_rom(2517)),16);
when x"9d6" => lut_sig <= to_unsigned(integer(my_rom(2518)),16);
when x"9d7" => lut_sig <= to_unsigned(integer(my_rom(2519)),16);
when x"9d8" => lut_sig <= to_unsigned(integer(my_rom(2520)),16);
when x"9d9" => lut_sig <= to_unsigned(integer(my_rom(2521)),16);
when x"9da" => lut_sig <= to_unsigned(integer(my_rom(2522)),16);
when x"9db" => lut_sig <= to_unsigned(integer(my_rom(2523)),16);
when x"9dc" => lut_sig <= to_unsigned(integer(my_rom(2524)),16);
when x"9dd" => lut_sig <= to_unsigned(integer(my_rom(2525)),16);
when x"9de" => lut_sig <= to_unsigned(integer(my_rom(2526)),16);
when x"9df" => lut_sig <= to_unsigned(integer(my_rom(2527)),16);
when x"9e0" => lut_sig <= to_unsigned(integer(my_rom(2528)),16);
when x"9e1" => lut_sig <= to_unsigned(integer(my_rom(2529)),16);
when x"9e2" => lut_sig <= to_unsigned(integer(my_rom(2530)),16);
when x"9e3" => lut_sig <= to_unsigned(integer(my_rom(2531)),16);
when x"9e4" => lut_sig <= to_unsigned(integer(my_rom(2532)),16);
when x"9e5" => lut_sig <= to_unsigned(integer(my_rom(2533)),16);
when x"9e6" => lut_sig <= to_unsigned(integer(my_rom(2534)),16);
when x"9e7" => lut_sig <= to_unsigned(integer(my_rom(2535)),16);
when x"9e8" => lut_sig <= to_unsigned(integer(my_rom(2536)),16);
when x"9e9" => lut_sig <= to_unsigned(integer(my_rom(2537)),16);
when x"9ea" => lut_sig <= to_unsigned(integer(my_rom(2538)),16);
when x"9eb" => lut_sig <= to_unsigned(integer(my_rom(2539)),16);
when x"9ec" => lut_sig <= to_unsigned(integer(my_rom(2540)),16);
when x"9ed" => lut_sig <= to_unsigned(integer(my_rom(2541)),16);
when x"9ee" => lut_sig <= to_unsigned(integer(my_rom(2542)),16);
when x"9ef" => lut_sig <= to_unsigned(integer(my_rom(2543)),16);
when x"9f0" => lut_sig <= to_unsigned(integer(my_rom(2544)),16);
when x"9f1" => lut_sig <= to_unsigned(integer(my_rom(2545)),16);
when x"9f2" => lut_sig <= to_unsigned(integer(my_rom(2546)),16);
when x"9f3" => lut_sig <= to_unsigned(integer(my_rom(2547)),16);
when x"9f4" => lut_sig <= to_unsigned(integer(my_rom(2548)),16);
when x"9f5" => lut_sig <= to_unsigned(integer(my_rom(2549)),16);
when x"9f6" => lut_sig <= to_unsigned(integer(my_rom(2550)),16);
when x"9f7" => lut_sig <= to_unsigned(integer(my_rom(2551)),16);
when x"9f8" => lut_sig <= to_unsigned(integer(my_rom(2552)),16);
when x"9f9" => lut_sig <= to_unsigned(integer(my_rom(2553)),16);
when x"9fa" => lut_sig <= to_unsigned(integer(my_rom(2554)),16);
when x"9fb" => lut_sig <= to_unsigned(integer(my_rom(2555)),16);
when x"9fc" => lut_sig <= to_unsigned(integer(my_rom(2556)),16);
when x"9fd" => lut_sig <= to_unsigned(integer(my_rom(2557)),16);
when x"9fe" => lut_sig <= to_unsigned(integer(my_rom(2558)),16);
when x"9ff" => lut_sig <= to_unsigned(integer(my_rom(2559)),16);
when x"a00" => lut_sig <= to_unsigned(integer(my_rom(2560)),16);
when x"a01" => lut_sig <= to_unsigned(integer(my_rom(2561)),16);
when x"a02" => lut_sig <= to_unsigned(integer(my_rom(2562)),16);
when x"a03" => lut_sig <= to_unsigned(integer(my_rom(2563)),16);
when x"a04" => lut_sig <= to_unsigned(integer(my_rom(2564)),16);
when x"a05" => lut_sig <= to_unsigned(integer(my_rom(2565)),16);
when x"a06" => lut_sig <= to_unsigned(integer(my_rom(2566)),16);
when x"a07" => lut_sig <= to_unsigned(integer(my_rom(2567)),16);
when x"a08" => lut_sig <= to_unsigned(integer(my_rom(2568)),16);
when x"a09" => lut_sig <= to_unsigned(integer(my_rom(2569)),16);
when x"a0a" => lut_sig <= to_unsigned(integer(my_rom(2570)),16);
when x"a0b" => lut_sig <= to_unsigned(integer(my_rom(2571)),16);
when x"a0c" => lut_sig <= to_unsigned(integer(my_rom(2572)),16);
when x"a0d" => lut_sig <= to_unsigned(integer(my_rom(2573)),16);
when x"a0e" => lut_sig <= to_unsigned(integer(my_rom(2574)),16);
when x"a0f" => lut_sig <= to_unsigned(integer(my_rom(2575)),16);
when x"a10" => lut_sig <= to_unsigned(integer(my_rom(2576)),16);
when x"a11" => lut_sig <= to_unsigned(integer(my_rom(2577)),16);
when x"a12" => lut_sig <= to_unsigned(integer(my_rom(2578)),16);
when x"a13" => lut_sig <= to_unsigned(integer(my_rom(2579)),16);
when x"a14" => lut_sig <= to_unsigned(integer(my_rom(2580)),16);
when x"a15" => lut_sig <= to_unsigned(integer(my_rom(2581)),16);
when x"a16" => lut_sig <= to_unsigned(integer(my_rom(2582)),16);
when x"a17" => lut_sig <= to_unsigned(integer(my_rom(2583)),16);
when x"a18" => lut_sig <= to_unsigned(integer(my_rom(2584)),16);
when x"a19" => lut_sig <= to_unsigned(integer(my_rom(2585)),16);
when x"a1a" => lut_sig <= to_unsigned(integer(my_rom(2586)),16);
when x"a1b" => lut_sig <= to_unsigned(integer(my_rom(2587)),16);
when x"a1c" => lut_sig <= to_unsigned(integer(my_rom(2588)),16);
when x"a1d" => lut_sig <= to_unsigned(integer(my_rom(2589)),16);
when x"a1e" => lut_sig <= to_unsigned(integer(my_rom(2590)),16);
when x"a1f" => lut_sig <= to_unsigned(integer(my_rom(2591)),16);
when x"a20" => lut_sig <= to_unsigned(integer(my_rom(2592)),16);
when x"a21" => lut_sig <= to_unsigned(integer(my_rom(2593)),16);
when x"a22" => lut_sig <= to_unsigned(integer(my_rom(2594)),16);
when x"a23" => lut_sig <= to_unsigned(integer(my_rom(2595)),16);
when x"a24" => lut_sig <= to_unsigned(integer(my_rom(2596)),16);
when x"a25" => lut_sig <= to_unsigned(integer(my_rom(2597)),16);
when x"a26" => lut_sig <= to_unsigned(integer(my_rom(2598)),16);
when x"a27" => lut_sig <= to_unsigned(integer(my_rom(2599)),16);
when x"a28" => lut_sig <= to_unsigned(integer(my_rom(2600)),16);
when x"a29" => lut_sig <= to_unsigned(integer(my_rom(2601)),16);
when x"a2a" => lut_sig <= to_unsigned(integer(my_rom(2602)),16);
when x"a2b" => lut_sig <= to_unsigned(integer(my_rom(2603)),16);
when x"a2c" => lut_sig <= to_unsigned(integer(my_rom(2604)),16);
when x"a2d" => lut_sig <= to_unsigned(integer(my_rom(2605)),16);
when x"a2e" => lut_sig <= to_unsigned(integer(my_rom(2606)),16);
when x"a2f" => lut_sig <= to_unsigned(integer(my_rom(2607)),16);
when x"a30" => lut_sig <= to_unsigned(integer(my_rom(2608)),16);
when x"a31" => lut_sig <= to_unsigned(integer(my_rom(2609)),16);
when x"a32" => lut_sig <= to_unsigned(integer(my_rom(2610)),16);
when x"a33" => lut_sig <= to_unsigned(integer(my_rom(2611)),16);
when x"a34" => lut_sig <= to_unsigned(integer(my_rom(2612)),16);
when x"a35" => lut_sig <= to_unsigned(integer(my_rom(2613)),16);
when x"a36" => lut_sig <= to_unsigned(integer(my_rom(2614)),16);
when x"a37" => lut_sig <= to_unsigned(integer(my_rom(2615)),16);
when x"a38" => lut_sig <= to_unsigned(integer(my_rom(2616)),16);
when x"a39" => lut_sig <= to_unsigned(integer(my_rom(2617)),16);
when x"a3a" => lut_sig <= to_unsigned(integer(my_rom(2618)),16);
when x"a3b" => lut_sig <= to_unsigned(integer(my_rom(2619)),16);
when x"a3c" => lut_sig <= to_unsigned(integer(my_rom(2620)),16);
when x"a3d" => lut_sig <= to_unsigned(integer(my_rom(2621)),16);
when x"a3e" => lut_sig <= to_unsigned(integer(my_rom(2622)),16);
when x"a3f" => lut_sig <= to_unsigned(integer(my_rom(2623)),16);
when x"a40" => lut_sig <= to_unsigned(integer(my_rom(2624)),16);
when x"a41" => lut_sig <= to_unsigned(integer(my_rom(2625)),16);
when x"a42" => lut_sig <= to_unsigned(integer(my_rom(2626)),16);
when x"a43" => lut_sig <= to_unsigned(integer(my_rom(2627)),16);
when x"a44" => lut_sig <= to_unsigned(integer(my_rom(2628)),16);
when x"a45" => lut_sig <= to_unsigned(integer(my_rom(2629)),16);
when x"a46" => lut_sig <= to_unsigned(integer(my_rom(2630)),16);
when x"a47" => lut_sig <= to_unsigned(integer(my_rom(2631)),16);
when x"a48" => lut_sig <= to_unsigned(integer(my_rom(2632)),16);
when x"a49" => lut_sig <= to_unsigned(integer(my_rom(2633)),16);
when x"a4a" => lut_sig <= to_unsigned(integer(my_rom(2634)),16);
when x"a4b" => lut_sig <= to_unsigned(integer(my_rom(2635)),16);
when x"a4c" => lut_sig <= to_unsigned(integer(my_rom(2636)),16);
when x"a4d" => lut_sig <= to_unsigned(integer(my_rom(2637)),16);
when x"a4e" => lut_sig <= to_unsigned(integer(my_rom(2638)),16);
when x"a4f" => lut_sig <= to_unsigned(integer(my_rom(2639)),16);
when x"a50" => lut_sig <= to_unsigned(integer(my_rom(2640)),16);
when x"a51" => lut_sig <= to_unsigned(integer(my_rom(2641)),16);
when x"a52" => lut_sig <= to_unsigned(integer(my_rom(2642)),16);
when x"a53" => lut_sig <= to_unsigned(integer(my_rom(2643)),16);
when x"a54" => lut_sig <= to_unsigned(integer(my_rom(2644)),16);
when x"a55" => lut_sig <= to_unsigned(integer(my_rom(2645)),16);
when x"a56" => lut_sig <= to_unsigned(integer(my_rom(2646)),16);
when x"a57" => lut_sig <= to_unsigned(integer(my_rom(2647)),16);
when x"a58" => lut_sig <= to_unsigned(integer(my_rom(2648)),16);
when x"a59" => lut_sig <= to_unsigned(integer(my_rom(2649)),16);
when x"a5a" => lut_sig <= to_unsigned(integer(my_rom(2650)),16);
when x"a5b" => lut_sig <= to_unsigned(integer(my_rom(2651)),16);
when x"a5c" => lut_sig <= to_unsigned(integer(my_rom(2652)),16);
when x"a5d" => lut_sig <= to_unsigned(integer(my_rom(2653)),16);
when x"a5e" => lut_sig <= to_unsigned(integer(my_rom(2654)),16);
when x"a5f" => lut_sig <= to_unsigned(integer(my_rom(2655)),16);
when x"a60" => lut_sig <= to_unsigned(integer(my_rom(2656)),16);
when x"a61" => lut_sig <= to_unsigned(integer(my_rom(2657)),16);
when x"a62" => lut_sig <= to_unsigned(integer(my_rom(2658)),16);
when x"a63" => lut_sig <= to_unsigned(integer(my_rom(2659)),16);
when x"a64" => lut_sig <= to_unsigned(integer(my_rom(2660)),16);
when x"a65" => lut_sig <= to_unsigned(integer(my_rom(2661)),16);
when x"a66" => lut_sig <= to_unsigned(integer(my_rom(2662)),16);
when x"a67" => lut_sig <= to_unsigned(integer(my_rom(2663)),16);
when x"a68" => lut_sig <= to_unsigned(integer(my_rom(2664)),16);
when x"a69" => lut_sig <= to_unsigned(integer(my_rom(2665)),16);
when x"a6a" => lut_sig <= to_unsigned(integer(my_rom(2666)),16);
when x"a6b" => lut_sig <= to_unsigned(integer(my_rom(2667)),16);
when x"a6c" => lut_sig <= to_unsigned(integer(my_rom(2668)),16);
when x"a6d" => lut_sig <= to_unsigned(integer(my_rom(2669)),16);
when x"a6e" => lut_sig <= to_unsigned(integer(my_rom(2670)),16);
when x"a6f" => lut_sig <= to_unsigned(integer(my_rom(2671)),16);
when x"a70" => lut_sig <= to_unsigned(integer(my_rom(2672)),16);
when x"a71" => lut_sig <= to_unsigned(integer(my_rom(2673)),16);
when x"a72" => lut_sig <= to_unsigned(integer(my_rom(2674)),16);
when x"a73" => lut_sig <= to_unsigned(integer(my_rom(2675)),16);
when x"a74" => lut_sig <= to_unsigned(integer(my_rom(2676)),16);
when x"a75" => lut_sig <= to_unsigned(integer(my_rom(2677)),16);
when x"a76" => lut_sig <= to_unsigned(integer(my_rom(2678)),16);
when x"a77" => lut_sig <= to_unsigned(integer(my_rom(2679)),16);
when x"a78" => lut_sig <= to_unsigned(integer(my_rom(2680)),16);
when x"a79" => lut_sig <= to_unsigned(integer(my_rom(2681)),16);
when x"a7a" => lut_sig <= to_unsigned(integer(my_rom(2682)),16);
when x"a7b" => lut_sig <= to_unsigned(integer(my_rom(2683)),16);
when x"a7c" => lut_sig <= to_unsigned(integer(my_rom(2684)),16);
when x"a7d" => lut_sig <= to_unsigned(integer(my_rom(2685)),16);
when x"a7e" => lut_sig <= to_unsigned(integer(my_rom(2686)),16);
when x"a7f" => lut_sig <= to_unsigned(integer(my_rom(2687)),16);
when x"a80" => lut_sig <= to_unsigned(integer(my_rom(2688)),16);
when x"a81" => lut_sig <= to_unsigned(integer(my_rom(2689)),16);
when x"a82" => lut_sig <= to_unsigned(integer(my_rom(2690)),16);
when x"a83" => lut_sig <= to_unsigned(integer(my_rom(2691)),16);
when x"a84" => lut_sig <= to_unsigned(integer(my_rom(2692)),16);
when x"a85" => lut_sig <= to_unsigned(integer(my_rom(2693)),16);
when x"a86" => lut_sig <= to_unsigned(integer(my_rom(2694)),16);
when x"a87" => lut_sig <= to_unsigned(integer(my_rom(2695)),16);
when x"a88" => lut_sig <= to_unsigned(integer(my_rom(2696)),16);
when x"a89" => lut_sig <= to_unsigned(integer(my_rom(2697)),16);
when x"a8a" => lut_sig <= to_unsigned(integer(my_rom(2698)),16);
when x"a8b" => lut_sig <= to_unsigned(integer(my_rom(2699)),16);
when x"a8c" => lut_sig <= to_unsigned(integer(my_rom(2700)),16);
when x"a8d" => lut_sig <= to_unsigned(integer(my_rom(2701)),16);
when x"a8e" => lut_sig <= to_unsigned(integer(my_rom(2702)),16);
when x"a8f" => lut_sig <= to_unsigned(integer(my_rom(2703)),16);
when x"a90" => lut_sig <= to_unsigned(integer(my_rom(2704)),16);
when x"a91" => lut_sig <= to_unsigned(integer(my_rom(2705)),16);
when x"a92" => lut_sig <= to_unsigned(integer(my_rom(2706)),16);
when x"a93" => lut_sig <= to_unsigned(integer(my_rom(2707)),16);
when x"a94" => lut_sig <= to_unsigned(integer(my_rom(2708)),16);
when x"a95" => lut_sig <= to_unsigned(integer(my_rom(2709)),16);
when x"a96" => lut_sig <= to_unsigned(integer(my_rom(2710)),16);
when x"a97" => lut_sig <= to_unsigned(integer(my_rom(2711)),16);
when x"a98" => lut_sig <= to_unsigned(integer(my_rom(2712)),16);
when x"a99" => lut_sig <= to_unsigned(integer(my_rom(2713)),16);
when x"a9a" => lut_sig <= to_unsigned(integer(my_rom(2714)),16);
when x"a9b" => lut_sig <= to_unsigned(integer(my_rom(2715)),16);
when x"a9c" => lut_sig <= to_unsigned(integer(my_rom(2716)),16);
when x"a9d" => lut_sig <= to_unsigned(integer(my_rom(2717)),16);
when x"a9e" => lut_sig <= to_unsigned(integer(my_rom(2718)),16);
when x"a9f" => lut_sig <= to_unsigned(integer(my_rom(2719)),16);
when x"aa0" => lut_sig <= to_unsigned(integer(my_rom(2720)),16);
when x"aa1" => lut_sig <= to_unsigned(integer(my_rom(2721)),16);
when x"aa2" => lut_sig <= to_unsigned(integer(my_rom(2722)),16);
when x"aa3" => lut_sig <= to_unsigned(integer(my_rom(2723)),16);
when x"aa4" => lut_sig <= to_unsigned(integer(my_rom(2724)),16);
when x"aa5" => lut_sig <= to_unsigned(integer(my_rom(2725)),16);
when x"aa6" => lut_sig <= to_unsigned(integer(my_rom(2726)),16);
when x"aa7" => lut_sig <= to_unsigned(integer(my_rom(2727)),16);
when x"aa8" => lut_sig <= to_unsigned(integer(my_rom(2728)),16);
when x"aa9" => lut_sig <= to_unsigned(integer(my_rom(2729)),16);
when x"aaa" => lut_sig <= to_unsigned(integer(my_rom(2730)),16);
when x"aab" => lut_sig <= to_unsigned(integer(my_rom(2731)),16);
when x"aac" => lut_sig <= to_unsigned(integer(my_rom(2732)),16);
when x"aad" => lut_sig <= to_unsigned(integer(my_rom(2733)),16);
when x"aae" => lut_sig <= to_unsigned(integer(my_rom(2734)),16);
when x"aaf" => lut_sig <= to_unsigned(integer(my_rom(2735)),16);
when x"ab0" => lut_sig <= to_unsigned(integer(my_rom(2736)),16);
when x"ab1" => lut_sig <= to_unsigned(integer(my_rom(2737)),16);
when x"ab2" => lut_sig <= to_unsigned(integer(my_rom(2738)),16);
when x"ab3" => lut_sig <= to_unsigned(integer(my_rom(2739)),16);
when x"ab4" => lut_sig <= to_unsigned(integer(my_rom(2740)),16);
when x"ab5" => lut_sig <= to_unsigned(integer(my_rom(2741)),16);
when x"ab6" => lut_sig <= to_unsigned(integer(my_rom(2742)),16);
when x"ab7" => lut_sig <= to_unsigned(integer(my_rom(2743)),16);
when x"ab8" => lut_sig <= to_unsigned(integer(my_rom(2744)),16);
when x"ab9" => lut_sig <= to_unsigned(integer(my_rom(2745)),16);
when x"aba" => lut_sig <= to_unsigned(integer(my_rom(2746)),16);
when x"abb" => lut_sig <= to_unsigned(integer(my_rom(2747)),16);
when x"abc" => lut_sig <= to_unsigned(integer(my_rom(2748)),16);
when x"abd" => lut_sig <= to_unsigned(integer(my_rom(2749)),16);
when x"abe" => lut_sig <= to_unsigned(integer(my_rom(2750)),16);
when x"abf" => lut_sig <= to_unsigned(integer(my_rom(2751)),16);
when x"ac0" => lut_sig <= to_unsigned(integer(my_rom(2752)),16);
when x"ac1" => lut_sig <= to_unsigned(integer(my_rom(2753)),16);
when x"ac2" => lut_sig <= to_unsigned(integer(my_rom(2754)),16);
when x"ac3" => lut_sig <= to_unsigned(integer(my_rom(2755)),16);
when x"ac4" => lut_sig <= to_unsigned(integer(my_rom(2756)),16);
when x"ac5" => lut_sig <= to_unsigned(integer(my_rom(2757)),16);
when x"ac6" => lut_sig <= to_unsigned(integer(my_rom(2758)),16);
when x"ac7" => lut_sig <= to_unsigned(integer(my_rom(2759)),16);
when x"ac8" => lut_sig <= to_unsigned(integer(my_rom(2760)),16);
when x"ac9" => lut_sig <= to_unsigned(integer(my_rom(2761)),16);
when x"aca" => lut_sig <= to_unsigned(integer(my_rom(2762)),16);
when x"acb" => lut_sig <= to_unsigned(integer(my_rom(2763)),16);
when x"acc" => lut_sig <= to_unsigned(integer(my_rom(2764)),16);
when x"acd" => lut_sig <= to_unsigned(integer(my_rom(2765)),16);
when x"ace" => lut_sig <= to_unsigned(integer(my_rom(2766)),16);
when x"acf" => lut_sig <= to_unsigned(integer(my_rom(2767)),16);
when x"ad0" => lut_sig <= to_unsigned(integer(my_rom(2768)),16);
when x"ad1" => lut_sig <= to_unsigned(integer(my_rom(2769)),16);
when x"ad2" => lut_sig <= to_unsigned(integer(my_rom(2770)),16);
when x"ad3" => lut_sig <= to_unsigned(integer(my_rom(2771)),16);
when x"ad4" => lut_sig <= to_unsigned(integer(my_rom(2772)),16);
when x"ad5" => lut_sig <= to_unsigned(integer(my_rom(2773)),16);
when x"ad6" => lut_sig <= to_unsigned(integer(my_rom(2774)),16);
when x"ad7" => lut_sig <= to_unsigned(integer(my_rom(2775)),16);
when x"ad8" => lut_sig <= to_unsigned(integer(my_rom(2776)),16);
when x"ad9" => lut_sig <= to_unsigned(integer(my_rom(2777)),16);
when x"ada" => lut_sig <= to_unsigned(integer(my_rom(2778)),16);
when x"adb" => lut_sig <= to_unsigned(integer(my_rom(2779)),16);
when x"adc" => lut_sig <= to_unsigned(integer(my_rom(2780)),16);
when x"add" => lut_sig <= to_unsigned(integer(my_rom(2781)),16);
when x"ade" => lut_sig <= to_unsigned(integer(my_rom(2782)),16);
when x"adf" => lut_sig <= to_unsigned(integer(my_rom(2783)),16);
when x"ae0" => lut_sig <= to_unsigned(integer(my_rom(2784)),16);
when x"ae1" => lut_sig <= to_unsigned(integer(my_rom(2785)),16);
when x"ae2" => lut_sig <= to_unsigned(integer(my_rom(2786)),16);
when x"ae3" => lut_sig <= to_unsigned(integer(my_rom(2787)),16);
when x"ae4" => lut_sig <= to_unsigned(integer(my_rom(2788)),16);
when x"ae5" => lut_sig <= to_unsigned(integer(my_rom(2789)),16);
when x"ae6" => lut_sig <= to_unsigned(integer(my_rom(2790)),16);
when x"ae7" => lut_sig <= to_unsigned(integer(my_rom(2791)),16);
when x"ae8" => lut_sig <= to_unsigned(integer(my_rom(2792)),16);
when x"ae9" => lut_sig <= to_unsigned(integer(my_rom(2793)),16);
when x"aea" => lut_sig <= to_unsigned(integer(my_rom(2794)),16);
when x"aeb" => lut_sig <= to_unsigned(integer(my_rom(2795)),16);
when x"aec" => lut_sig <= to_unsigned(integer(my_rom(2796)),16);
when x"aed" => lut_sig <= to_unsigned(integer(my_rom(2797)),16);
when x"aee" => lut_sig <= to_unsigned(integer(my_rom(2798)),16);
when x"aef" => lut_sig <= to_unsigned(integer(my_rom(2799)),16);
when x"af0" => lut_sig <= to_unsigned(integer(my_rom(2800)),16);
when x"af1" => lut_sig <= to_unsigned(integer(my_rom(2801)),16);
when x"af2" => lut_sig <= to_unsigned(integer(my_rom(2802)),16);
when x"af3" => lut_sig <= to_unsigned(integer(my_rom(2803)),16);
when x"af4" => lut_sig <= to_unsigned(integer(my_rom(2804)),16);
when x"af5" => lut_sig <= to_unsigned(integer(my_rom(2805)),16);
when x"af6" => lut_sig <= to_unsigned(integer(my_rom(2806)),16);
when x"af7" => lut_sig <= to_unsigned(integer(my_rom(2807)),16);
when x"af8" => lut_sig <= to_unsigned(integer(my_rom(2808)),16);
when x"af9" => lut_sig <= to_unsigned(integer(my_rom(2809)),16);
when x"afa" => lut_sig <= to_unsigned(integer(my_rom(2810)),16);
when x"afb" => lut_sig <= to_unsigned(integer(my_rom(2811)),16);
when x"afc" => lut_sig <= to_unsigned(integer(my_rom(2812)),16);
when x"afd" => lut_sig <= to_unsigned(integer(my_rom(2813)),16);
when x"afe" => lut_sig <= to_unsigned(integer(my_rom(2814)),16);
when x"aff" => lut_sig <= to_unsigned(integer(my_rom(2815)),16);
when x"b00" => lut_sig <= to_unsigned(integer(my_rom(2816)),16);
when x"b01" => lut_sig <= to_unsigned(integer(my_rom(2817)),16);
when x"b02" => lut_sig <= to_unsigned(integer(my_rom(2818)),16);
when x"b03" => lut_sig <= to_unsigned(integer(my_rom(2819)),16);
when x"b04" => lut_sig <= to_unsigned(integer(my_rom(2820)),16);
when x"b05" => lut_sig <= to_unsigned(integer(my_rom(2821)),16);
when x"b06" => lut_sig <= to_unsigned(integer(my_rom(2822)),16);
when x"b07" => lut_sig <= to_unsigned(integer(my_rom(2823)),16);
when x"b08" => lut_sig <= to_unsigned(integer(my_rom(2824)),16);
when x"b09" => lut_sig <= to_unsigned(integer(my_rom(2825)),16);
when x"b0a" => lut_sig <= to_unsigned(integer(my_rom(2826)),16);
when x"b0b" => lut_sig <= to_unsigned(integer(my_rom(2827)),16);
when x"b0c" => lut_sig <= to_unsigned(integer(my_rom(2828)),16);
when x"b0d" => lut_sig <= to_unsigned(integer(my_rom(2829)),16);
when x"b0e" => lut_sig <= to_unsigned(integer(my_rom(2830)),16);
when x"b0f" => lut_sig <= to_unsigned(integer(my_rom(2831)),16);
when x"b10" => lut_sig <= to_unsigned(integer(my_rom(2832)),16);
when x"b11" => lut_sig <= to_unsigned(integer(my_rom(2833)),16);
when x"b12" => lut_sig <= to_unsigned(integer(my_rom(2834)),16);
when x"b13" => lut_sig <= to_unsigned(integer(my_rom(2835)),16);
when x"b14" => lut_sig <= to_unsigned(integer(my_rom(2836)),16);
when x"b15" => lut_sig <= to_unsigned(integer(my_rom(2837)),16);
when x"b16" => lut_sig <= to_unsigned(integer(my_rom(2838)),16);
when x"b17" => lut_sig <= to_unsigned(integer(my_rom(2839)),16);
when x"b18" => lut_sig <= to_unsigned(integer(my_rom(2840)),16);
when x"b19" => lut_sig <= to_unsigned(integer(my_rom(2841)),16);
when x"b1a" => lut_sig <= to_unsigned(integer(my_rom(2842)),16);
when x"b1b" => lut_sig <= to_unsigned(integer(my_rom(2843)),16);
when x"b1c" => lut_sig <= to_unsigned(integer(my_rom(2844)),16);
when x"b1d" => lut_sig <= to_unsigned(integer(my_rom(2845)),16);
when x"b1e" => lut_sig <= to_unsigned(integer(my_rom(2846)),16);
when x"b1f" => lut_sig <= to_unsigned(integer(my_rom(2847)),16);
when x"b20" => lut_sig <= to_unsigned(integer(my_rom(2848)),16);
when x"b21" => lut_sig <= to_unsigned(integer(my_rom(2849)),16);
when x"b22" => lut_sig <= to_unsigned(integer(my_rom(2850)),16);
when x"b23" => lut_sig <= to_unsigned(integer(my_rom(2851)),16);
when x"b24" => lut_sig <= to_unsigned(integer(my_rom(2852)),16);
when x"b25" => lut_sig <= to_unsigned(integer(my_rom(2853)),16);
when x"b26" => lut_sig <= to_unsigned(integer(my_rom(2854)),16);
when x"b27" => lut_sig <= to_unsigned(integer(my_rom(2855)),16);
when x"b28" => lut_sig <= to_unsigned(integer(my_rom(2856)),16);
when x"b29" => lut_sig <= to_unsigned(integer(my_rom(2857)),16);
when x"b2a" => lut_sig <= to_unsigned(integer(my_rom(2858)),16);
when x"b2b" => lut_sig <= to_unsigned(integer(my_rom(2859)),16);
when x"b2c" => lut_sig <= to_unsigned(integer(my_rom(2860)),16);
when x"b2d" => lut_sig <= to_unsigned(integer(my_rom(2861)),16);
when x"b2e" => lut_sig <= to_unsigned(integer(my_rom(2862)),16);
when x"b2f" => lut_sig <= to_unsigned(integer(my_rom(2863)),16);
when x"b30" => lut_sig <= to_unsigned(integer(my_rom(2864)),16);
when x"b31" => lut_sig <= to_unsigned(integer(my_rom(2865)),16);
when x"b32" => lut_sig <= to_unsigned(integer(my_rom(2866)),16);
when x"b33" => lut_sig <= to_unsigned(integer(my_rom(2867)),16);
when x"b34" => lut_sig <= to_unsigned(integer(my_rom(2868)),16);
when x"b35" => lut_sig <= to_unsigned(integer(my_rom(2869)),16);
when x"b36" => lut_sig <= to_unsigned(integer(my_rom(2870)),16);
when x"b37" => lut_sig <= to_unsigned(integer(my_rom(2871)),16);
when x"b38" => lut_sig <= to_unsigned(integer(my_rom(2872)),16);
when x"b39" => lut_sig <= to_unsigned(integer(my_rom(2873)),16);
when x"b3a" => lut_sig <= to_unsigned(integer(my_rom(2874)),16);
when x"b3b" => lut_sig <= to_unsigned(integer(my_rom(2875)),16);
when x"b3c" => lut_sig <= to_unsigned(integer(my_rom(2876)),16);
when x"b3d" => lut_sig <= to_unsigned(integer(my_rom(2877)),16);
when x"b3e" => lut_sig <= to_unsigned(integer(my_rom(2878)),16);
when x"b3f" => lut_sig <= to_unsigned(integer(my_rom(2879)),16);
when x"b40" => lut_sig <= to_unsigned(integer(my_rom(2880)),16);
when x"b41" => lut_sig <= to_unsigned(integer(my_rom(2881)),16);
when x"b42" => lut_sig <= to_unsigned(integer(my_rom(2882)),16);
when x"b43" => lut_sig <= to_unsigned(integer(my_rom(2883)),16);
when x"b44" => lut_sig <= to_unsigned(integer(my_rom(2884)),16);
when x"b45" => lut_sig <= to_unsigned(integer(my_rom(2885)),16);
when x"b46" => lut_sig <= to_unsigned(integer(my_rom(2886)),16);
when x"b47" => lut_sig <= to_unsigned(integer(my_rom(2887)),16);
when x"b48" => lut_sig <= to_unsigned(integer(my_rom(2888)),16);
when x"b49" => lut_sig <= to_unsigned(integer(my_rom(2889)),16);
when x"b4a" => lut_sig <= to_unsigned(integer(my_rom(2890)),16);
when x"b4b" => lut_sig <= to_unsigned(integer(my_rom(2891)),16);
when x"b4c" => lut_sig <= to_unsigned(integer(my_rom(2892)),16);
when x"b4d" => lut_sig <= to_unsigned(integer(my_rom(2893)),16);
when x"b4e" => lut_sig <= to_unsigned(integer(my_rom(2894)),16);
when x"b4f" => lut_sig <= to_unsigned(integer(my_rom(2895)),16);
when x"b50" => lut_sig <= to_unsigned(integer(my_rom(2896)),16);
when x"b51" => lut_sig <= to_unsigned(integer(my_rom(2897)),16);
when x"b52" => lut_sig <= to_unsigned(integer(my_rom(2898)),16);
when x"b53" => lut_sig <= to_unsigned(integer(my_rom(2899)),16);
when x"b54" => lut_sig <= to_unsigned(integer(my_rom(2900)),16);
when x"b55" => lut_sig <= to_unsigned(integer(my_rom(2901)),16);
when x"b56" => lut_sig <= to_unsigned(integer(my_rom(2902)),16);
when x"b57" => lut_sig <= to_unsigned(integer(my_rom(2903)),16);
when x"b58" => lut_sig <= to_unsigned(integer(my_rom(2904)),16);
when x"b59" => lut_sig <= to_unsigned(integer(my_rom(2905)),16);
when x"b5a" => lut_sig <= to_unsigned(integer(my_rom(2906)),16);
when x"b5b" => lut_sig <= to_unsigned(integer(my_rom(2907)),16);
when x"b5c" => lut_sig <= to_unsigned(integer(my_rom(2908)),16);
when x"b5d" => lut_sig <= to_unsigned(integer(my_rom(2909)),16);
when x"b5e" => lut_sig <= to_unsigned(integer(my_rom(2910)),16);
when x"b5f" => lut_sig <= to_unsigned(integer(my_rom(2911)),16);
when x"b60" => lut_sig <= to_unsigned(integer(my_rom(2912)),16);
when x"b61" => lut_sig <= to_unsigned(integer(my_rom(2913)),16);
when x"b62" => lut_sig <= to_unsigned(integer(my_rom(2914)),16);
when x"b63" => lut_sig <= to_unsigned(integer(my_rom(2915)),16);
when x"b64" => lut_sig <= to_unsigned(integer(my_rom(2916)),16);
when x"b65" => lut_sig <= to_unsigned(integer(my_rom(2917)),16);
when x"b66" => lut_sig <= to_unsigned(integer(my_rom(2918)),16);
when x"b67" => lut_sig <= to_unsigned(integer(my_rom(2919)),16);
when x"b68" => lut_sig <= to_unsigned(integer(my_rom(2920)),16);
when x"b69" => lut_sig <= to_unsigned(integer(my_rom(2921)),16);
when x"b6a" => lut_sig <= to_unsigned(integer(my_rom(2922)),16);
when x"b6b" => lut_sig <= to_unsigned(integer(my_rom(2923)),16);
when x"b6c" => lut_sig <= to_unsigned(integer(my_rom(2924)),16);
when x"b6d" => lut_sig <= to_unsigned(integer(my_rom(2925)),16);
when x"b6e" => lut_sig <= to_unsigned(integer(my_rom(2926)),16);
when x"b6f" => lut_sig <= to_unsigned(integer(my_rom(2927)),16);
when x"b70" => lut_sig <= to_unsigned(integer(my_rom(2928)),16);
when x"b71" => lut_sig <= to_unsigned(integer(my_rom(2929)),16);
when x"b72" => lut_sig <= to_unsigned(integer(my_rom(2930)),16);
when x"b73" => lut_sig <= to_unsigned(integer(my_rom(2931)),16);
when x"b74" => lut_sig <= to_unsigned(integer(my_rom(2932)),16);
when x"b75" => lut_sig <= to_unsigned(integer(my_rom(2933)),16);
when x"b76" => lut_sig <= to_unsigned(integer(my_rom(2934)),16);
when x"b77" => lut_sig <= to_unsigned(integer(my_rom(2935)),16);
when x"b78" => lut_sig <= to_unsigned(integer(my_rom(2936)),16);
when x"b79" => lut_sig <= to_unsigned(integer(my_rom(2937)),16);
when x"b7a" => lut_sig <= to_unsigned(integer(my_rom(2938)),16);
when x"b7b" => lut_sig <= to_unsigned(integer(my_rom(2939)),16);
when x"b7c" => lut_sig <= to_unsigned(integer(my_rom(2940)),16);
when x"b7d" => lut_sig <= to_unsigned(integer(my_rom(2941)),16);
when x"b7e" => lut_sig <= to_unsigned(integer(my_rom(2942)),16);
when x"b7f" => lut_sig <= to_unsigned(integer(my_rom(2943)),16);
when x"b80" => lut_sig <= to_unsigned(integer(my_rom(2944)),16);
when x"b81" => lut_sig <= to_unsigned(integer(my_rom(2945)),16);
when x"b82" => lut_sig <= to_unsigned(integer(my_rom(2946)),16);
when x"b83" => lut_sig <= to_unsigned(integer(my_rom(2947)),16);
when x"b84" => lut_sig <= to_unsigned(integer(my_rom(2948)),16);
when x"b85" => lut_sig <= to_unsigned(integer(my_rom(2949)),16);
when x"b86" => lut_sig <= to_unsigned(integer(my_rom(2950)),16);
when x"b87" => lut_sig <= to_unsigned(integer(my_rom(2951)),16);
when x"b88" => lut_sig <= to_unsigned(integer(my_rom(2952)),16);
when x"b89" => lut_sig <= to_unsigned(integer(my_rom(2953)),16);
when x"b8a" => lut_sig <= to_unsigned(integer(my_rom(2954)),16);
when x"b8b" => lut_sig <= to_unsigned(integer(my_rom(2955)),16);
when x"b8c" => lut_sig <= to_unsigned(integer(my_rom(2956)),16);
when x"b8d" => lut_sig <= to_unsigned(integer(my_rom(2957)),16);
when x"b8e" => lut_sig <= to_unsigned(integer(my_rom(2958)),16);
when x"b8f" => lut_sig <= to_unsigned(integer(my_rom(2959)),16);
when x"b90" => lut_sig <= to_unsigned(integer(my_rom(2960)),16);
when x"b91" => lut_sig <= to_unsigned(integer(my_rom(2961)),16);
when x"b92" => lut_sig <= to_unsigned(integer(my_rom(2962)),16);
when x"b93" => lut_sig <= to_unsigned(integer(my_rom(2963)),16);
when x"b94" => lut_sig <= to_unsigned(integer(my_rom(2964)),16);
when x"b95" => lut_sig <= to_unsigned(integer(my_rom(2965)),16);
when x"b96" => lut_sig <= to_unsigned(integer(my_rom(2966)),16);
when x"b97" => lut_sig <= to_unsigned(integer(my_rom(2967)),16);
when x"b98" => lut_sig <= to_unsigned(integer(my_rom(2968)),16);
when x"b99" => lut_sig <= to_unsigned(integer(my_rom(2969)),16);
when x"b9a" => lut_sig <= to_unsigned(integer(my_rom(2970)),16);
when x"b9b" => lut_sig <= to_unsigned(integer(my_rom(2971)),16);
when x"b9c" => lut_sig <= to_unsigned(integer(my_rom(2972)),16);
when x"b9d" => lut_sig <= to_unsigned(integer(my_rom(2973)),16);
when x"b9e" => lut_sig <= to_unsigned(integer(my_rom(2974)),16);
when x"b9f" => lut_sig <= to_unsigned(integer(my_rom(2975)),16);
when x"ba0" => lut_sig <= to_unsigned(integer(my_rom(2976)),16);
when x"ba1" => lut_sig <= to_unsigned(integer(my_rom(2977)),16);
when x"ba2" => lut_sig <= to_unsigned(integer(my_rom(2978)),16);
when x"ba3" => lut_sig <= to_unsigned(integer(my_rom(2979)),16);
when x"ba4" => lut_sig <= to_unsigned(integer(my_rom(2980)),16);
when x"ba5" => lut_sig <= to_unsigned(integer(my_rom(2981)),16);
when x"ba6" => lut_sig <= to_unsigned(integer(my_rom(2982)),16);
when x"ba7" => lut_sig <= to_unsigned(integer(my_rom(2983)),16);
when x"ba8" => lut_sig <= to_unsigned(integer(my_rom(2984)),16);
when x"ba9" => lut_sig <= to_unsigned(integer(my_rom(2985)),16);
when x"baa" => lut_sig <= to_unsigned(integer(my_rom(2986)),16);
when x"bab" => lut_sig <= to_unsigned(integer(my_rom(2987)),16);
when x"bac" => lut_sig <= to_unsigned(integer(my_rom(2988)),16);
when x"bad" => lut_sig <= to_unsigned(integer(my_rom(2989)),16);
when x"bae" => lut_sig <= to_unsigned(integer(my_rom(2990)),16);
when x"baf" => lut_sig <= to_unsigned(integer(my_rom(2991)),16);
when x"bb0" => lut_sig <= to_unsigned(integer(my_rom(2992)),16);
when x"bb1" => lut_sig <= to_unsigned(integer(my_rom(2993)),16);
when x"bb2" => lut_sig <= to_unsigned(integer(my_rom(2994)),16);
when x"bb3" => lut_sig <= to_unsigned(integer(my_rom(2995)),16);
when x"bb4" => lut_sig <= to_unsigned(integer(my_rom(2996)),16);
when x"bb5" => lut_sig <= to_unsigned(integer(my_rom(2997)),16);
when x"bb6" => lut_sig <= to_unsigned(integer(my_rom(2998)),16);
when x"bb7" => lut_sig <= to_unsigned(integer(my_rom(2999)),16);
when x"bb8" => lut_sig <= to_unsigned(integer(my_rom(3000)),16);
when x"bb9" => lut_sig <= to_unsigned(integer(my_rom(3001)),16);
when x"bba" => lut_sig <= to_unsigned(integer(my_rom(3002)),16);
when x"bbb" => lut_sig <= to_unsigned(integer(my_rom(3003)),16);
when x"bbc" => lut_sig <= to_unsigned(integer(my_rom(3004)),16);
when x"bbd" => lut_sig <= to_unsigned(integer(my_rom(3005)),16);
when x"bbe" => lut_sig <= to_unsigned(integer(my_rom(3006)),16);
when x"bbf" => lut_sig <= to_unsigned(integer(my_rom(3007)),16);
when x"bc0" => lut_sig <= to_unsigned(integer(my_rom(3008)),16);
when x"bc1" => lut_sig <= to_unsigned(integer(my_rom(3009)),16);
when x"bc2" => lut_sig <= to_unsigned(integer(my_rom(3010)),16);
when x"bc3" => lut_sig <= to_unsigned(integer(my_rom(3011)),16);
when x"bc4" => lut_sig <= to_unsigned(integer(my_rom(3012)),16);
when x"bc5" => lut_sig <= to_unsigned(integer(my_rom(3013)),16);
when x"bc6" => lut_sig <= to_unsigned(integer(my_rom(3014)),16);
when x"bc7" => lut_sig <= to_unsigned(integer(my_rom(3015)),16);
when x"bc8" => lut_sig <= to_unsigned(integer(my_rom(3016)),16);
when x"bc9" => lut_sig <= to_unsigned(integer(my_rom(3017)),16);
when x"bca" => lut_sig <= to_unsigned(integer(my_rom(3018)),16);
when x"bcb" => lut_sig <= to_unsigned(integer(my_rom(3019)),16);
when x"bcc" => lut_sig <= to_unsigned(integer(my_rom(3020)),16);
when x"bcd" => lut_sig <= to_unsigned(integer(my_rom(3021)),16);
when x"bce" => lut_sig <= to_unsigned(integer(my_rom(3022)),16);
when x"bcf" => lut_sig <= to_unsigned(integer(my_rom(3023)),16);
when x"bd0" => lut_sig <= to_unsigned(integer(my_rom(3024)),16);
when x"bd1" => lut_sig <= to_unsigned(integer(my_rom(3025)),16);
when x"bd2" => lut_sig <= to_unsigned(integer(my_rom(3026)),16);
when x"bd3" => lut_sig <= to_unsigned(integer(my_rom(3027)),16);
when x"bd4" => lut_sig <= to_unsigned(integer(my_rom(3028)),16);
when x"bd5" => lut_sig <= to_unsigned(integer(my_rom(3029)),16);
when x"bd6" => lut_sig <= to_unsigned(integer(my_rom(3030)),16);
when x"bd7" => lut_sig <= to_unsigned(integer(my_rom(3031)),16);
when x"bd8" => lut_sig <= to_unsigned(integer(my_rom(3032)),16);
when x"bd9" => lut_sig <= to_unsigned(integer(my_rom(3033)),16);
when x"bda" => lut_sig <= to_unsigned(integer(my_rom(3034)),16);
when x"bdb" => lut_sig <= to_unsigned(integer(my_rom(3035)),16);
when x"bdc" => lut_sig <= to_unsigned(integer(my_rom(3036)),16);
when x"bdd" => lut_sig <= to_unsigned(integer(my_rom(3037)),16);
when x"bde" => lut_sig <= to_unsigned(integer(my_rom(3038)),16);
when x"bdf" => lut_sig <= to_unsigned(integer(my_rom(3039)),16);
when x"be0" => lut_sig <= to_unsigned(integer(my_rom(3040)),16);
when x"be1" => lut_sig <= to_unsigned(integer(my_rom(3041)),16);
when x"be2" => lut_sig <= to_unsigned(integer(my_rom(3042)),16);
when x"be3" => lut_sig <= to_unsigned(integer(my_rom(3043)),16);
when x"be4" => lut_sig <= to_unsigned(integer(my_rom(3044)),16);
when x"be5" => lut_sig <= to_unsigned(integer(my_rom(3045)),16);
when x"be6" => lut_sig <= to_unsigned(integer(my_rom(3046)),16);
when x"be7" => lut_sig <= to_unsigned(integer(my_rom(3047)),16);
when x"be8" => lut_sig <= to_unsigned(integer(my_rom(3048)),16);
when x"be9" => lut_sig <= to_unsigned(integer(my_rom(3049)),16);
when x"bea" => lut_sig <= to_unsigned(integer(my_rom(3050)),16);
when x"beb" => lut_sig <= to_unsigned(integer(my_rom(3051)),16);
when x"bec" => lut_sig <= to_unsigned(integer(my_rom(3052)),16);
when x"bed" => lut_sig <= to_unsigned(integer(my_rom(3053)),16);
when x"bee" => lut_sig <= to_unsigned(integer(my_rom(3054)),16);
when x"bef" => lut_sig <= to_unsigned(integer(my_rom(3055)),16);
when x"bf0" => lut_sig <= to_unsigned(integer(my_rom(3056)),16);
when x"bf1" => lut_sig <= to_unsigned(integer(my_rom(3057)),16);
when x"bf2" => lut_sig <= to_unsigned(integer(my_rom(3058)),16);
when x"bf3" => lut_sig <= to_unsigned(integer(my_rom(3059)),16);
when x"bf4" => lut_sig <= to_unsigned(integer(my_rom(3060)),16);
when x"bf5" => lut_sig <= to_unsigned(integer(my_rom(3061)),16);
when x"bf6" => lut_sig <= to_unsigned(integer(my_rom(3062)),16);
when x"bf7" => lut_sig <= to_unsigned(integer(my_rom(3063)),16);
when x"bf8" => lut_sig <= to_unsigned(integer(my_rom(3064)),16);
when x"bf9" => lut_sig <= to_unsigned(integer(my_rom(3065)),16);
when x"bfa" => lut_sig <= to_unsigned(integer(my_rom(3066)),16);
when x"bfb" => lut_sig <= to_unsigned(integer(my_rom(3067)),16);
when x"bfc" => lut_sig <= to_unsigned(integer(my_rom(3068)),16);
when x"bfd" => lut_sig <= to_unsigned(integer(my_rom(3069)),16);
when x"bfe" => lut_sig <= to_unsigned(integer(my_rom(3070)),16);
when x"bff" => lut_sig <= to_unsigned(integer(my_rom(3071)),16);
when x"c00" => lut_sig <= to_unsigned(integer(my_rom(3072)),16);
when x"c01" => lut_sig <= to_unsigned(integer(my_rom(3073)),16);
when x"c02" => lut_sig <= to_unsigned(integer(my_rom(3074)),16);
when x"c03" => lut_sig <= to_unsigned(integer(my_rom(3075)),16);
when x"c04" => lut_sig <= to_unsigned(integer(my_rom(3076)),16);
when x"c05" => lut_sig <= to_unsigned(integer(my_rom(3077)),16);
when x"c06" => lut_sig <= to_unsigned(integer(my_rom(3078)),16);
when x"c07" => lut_sig <= to_unsigned(integer(my_rom(3079)),16);
when x"c08" => lut_sig <= to_unsigned(integer(my_rom(3080)),16);
when x"c09" => lut_sig <= to_unsigned(integer(my_rom(3081)),16);
when x"c0a" => lut_sig <= to_unsigned(integer(my_rom(3082)),16);
when x"c0b" => lut_sig <= to_unsigned(integer(my_rom(3083)),16);
when x"c0c" => lut_sig <= to_unsigned(integer(my_rom(3084)),16);
when x"c0d" => lut_sig <= to_unsigned(integer(my_rom(3085)),16);
when x"c0e" => lut_sig <= to_unsigned(integer(my_rom(3086)),16);
when x"c0f" => lut_sig <= to_unsigned(integer(my_rom(3087)),16);
when x"c10" => lut_sig <= to_unsigned(integer(my_rom(3088)),16);
when x"c11" => lut_sig <= to_unsigned(integer(my_rom(3089)),16);
when x"c12" => lut_sig <= to_unsigned(integer(my_rom(3090)),16);
when x"c13" => lut_sig <= to_unsigned(integer(my_rom(3091)),16);
when x"c14" => lut_sig <= to_unsigned(integer(my_rom(3092)),16);
when x"c15" => lut_sig <= to_unsigned(integer(my_rom(3093)),16);
when x"c16" => lut_sig <= to_unsigned(integer(my_rom(3094)),16);
when x"c17" => lut_sig <= to_unsigned(integer(my_rom(3095)),16);
when x"c18" => lut_sig <= to_unsigned(integer(my_rom(3096)),16);
when x"c19" => lut_sig <= to_unsigned(integer(my_rom(3097)),16);
when x"c1a" => lut_sig <= to_unsigned(integer(my_rom(3098)),16);
when x"c1b" => lut_sig <= to_unsigned(integer(my_rom(3099)),16);
when x"c1c" => lut_sig <= to_unsigned(integer(my_rom(3100)),16);
when x"c1d" => lut_sig <= to_unsigned(integer(my_rom(3101)),16);
when x"c1e" => lut_sig <= to_unsigned(integer(my_rom(3102)),16);
when x"c1f" => lut_sig <= to_unsigned(integer(my_rom(3103)),16);
when x"c20" => lut_sig <= to_unsigned(integer(my_rom(3104)),16);
when x"c21" => lut_sig <= to_unsigned(integer(my_rom(3105)),16);
when x"c22" => lut_sig <= to_unsigned(integer(my_rom(3106)),16);
when x"c23" => lut_sig <= to_unsigned(integer(my_rom(3107)),16);
when x"c24" => lut_sig <= to_unsigned(integer(my_rom(3108)),16);
when x"c25" => lut_sig <= to_unsigned(integer(my_rom(3109)),16);
when x"c26" => lut_sig <= to_unsigned(integer(my_rom(3110)),16);
when x"c27" => lut_sig <= to_unsigned(integer(my_rom(3111)),16);
when x"c28" => lut_sig <= to_unsigned(integer(my_rom(3112)),16);
when x"c29" => lut_sig <= to_unsigned(integer(my_rom(3113)),16);
when x"c2a" => lut_sig <= to_unsigned(integer(my_rom(3114)),16);
when x"c2b" => lut_sig <= to_unsigned(integer(my_rom(3115)),16);
when x"c2c" => lut_sig <= to_unsigned(integer(my_rom(3116)),16);
when x"c2d" => lut_sig <= to_unsigned(integer(my_rom(3117)),16);
when x"c2e" => lut_sig <= to_unsigned(integer(my_rom(3118)),16);
when x"c2f" => lut_sig <= to_unsigned(integer(my_rom(3119)),16);
when x"c30" => lut_sig <= to_unsigned(integer(my_rom(3120)),16);
when x"c31" => lut_sig <= to_unsigned(integer(my_rom(3121)),16);
when x"c32" => lut_sig <= to_unsigned(integer(my_rom(3122)),16);
when x"c33" => lut_sig <= to_unsigned(integer(my_rom(3123)),16);
when x"c34" => lut_sig <= to_unsigned(integer(my_rom(3124)),16);
when x"c35" => lut_sig <= to_unsigned(integer(my_rom(3125)),16);
when x"c36" => lut_sig <= to_unsigned(integer(my_rom(3126)),16);
when x"c37" => lut_sig <= to_unsigned(integer(my_rom(3127)),16);
when x"c38" => lut_sig <= to_unsigned(integer(my_rom(3128)),16);
when x"c39" => lut_sig <= to_unsigned(integer(my_rom(3129)),16);
when x"c3a" => lut_sig <= to_unsigned(integer(my_rom(3130)),16);
when x"c3b" => lut_sig <= to_unsigned(integer(my_rom(3131)),16);
when x"c3c" => lut_sig <= to_unsigned(integer(my_rom(3132)),16);
when x"c3d" => lut_sig <= to_unsigned(integer(my_rom(3133)),16);
when x"c3e" => lut_sig <= to_unsigned(integer(my_rom(3134)),16);
when x"c3f" => lut_sig <= to_unsigned(integer(my_rom(3135)),16);
when x"c40" => lut_sig <= to_unsigned(integer(my_rom(3136)),16);
when x"c41" => lut_sig <= to_unsigned(integer(my_rom(3137)),16);
when x"c42" => lut_sig <= to_unsigned(integer(my_rom(3138)),16);
when x"c43" => lut_sig <= to_unsigned(integer(my_rom(3139)),16);
when x"c44" => lut_sig <= to_unsigned(integer(my_rom(3140)),16);
when x"c45" => lut_sig <= to_unsigned(integer(my_rom(3141)),16);
when x"c46" => lut_sig <= to_unsigned(integer(my_rom(3142)),16);
when x"c47" => lut_sig <= to_unsigned(integer(my_rom(3143)),16);
when x"c48" => lut_sig <= to_unsigned(integer(my_rom(3144)),16);
when x"c49" => lut_sig <= to_unsigned(integer(my_rom(3145)),16);
when x"c4a" => lut_sig <= to_unsigned(integer(my_rom(3146)),16);
when x"c4b" => lut_sig <= to_unsigned(integer(my_rom(3147)),16);
when x"c4c" => lut_sig <= to_unsigned(integer(my_rom(3148)),16);
when x"c4d" => lut_sig <= to_unsigned(integer(my_rom(3149)),16);
when x"c4e" => lut_sig <= to_unsigned(integer(my_rom(3150)),16);
when x"c4f" => lut_sig <= to_unsigned(integer(my_rom(3151)),16);
when x"c50" => lut_sig <= to_unsigned(integer(my_rom(3152)),16);
when x"c51" => lut_sig <= to_unsigned(integer(my_rom(3153)),16);
when x"c52" => lut_sig <= to_unsigned(integer(my_rom(3154)),16);
when x"c53" => lut_sig <= to_unsigned(integer(my_rom(3155)),16);
when x"c54" => lut_sig <= to_unsigned(integer(my_rom(3156)),16);
when x"c55" => lut_sig <= to_unsigned(integer(my_rom(3157)),16);
when x"c56" => lut_sig <= to_unsigned(integer(my_rom(3158)),16);
when x"c57" => lut_sig <= to_unsigned(integer(my_rom(3159)),16);
when x"c58" => lut_sig <= to_unsigned(integer(my_rom(3160)),16);
when x"c59" => lut_sig <= to_unsigned(integer(my_rom(3161)),16);
when x"c5a" => lut_sig <= to_unsigned(integer(my_rom(3162)),16);
when x"c5b" => lut_sig <= to_unsigned(integer(my_rom(3163)),16);
when x"c5c" => lut_sig <= to_unsigned(integer(my_rom(3164)),16);
when x"c5d" => lut_sig <= to_unsigned(integer(my_rom(3165)),16);
when x"c5e" => lut_sig <= to_unsigned(integer(my_rom(3166)),16);
when x"c5f" => lut_sig <= to_unsigned(integer(my_rom(3167)),16);
when x"c60" => lut_sig <= to_unsigned(integer(my_rom(3168)),16);
when x"c61" => lut_sig <= to_unsigned(integer(my_rom(3169)),16);
when x"c62" => lut_sig <= to_unsigned(integer(my_rom(3170)),16);
when x"c63" => lut_sig <= to_unsigned(integer(my_rom(3171)),16);
when x"c64" => lut_sig <= to_unsigned(integer(my_rom(3172)),16);
when x"c65" => lut_sig <= to_unsigned(integer(my_rom(3173)),16);
when x"c66" => lut_sig <= to_unsigned(integer(my_rom(3174)),16);
when x"c67" => lut_sig <= to_unsigned(integer(my_rom(3175)),16);
when x"c68" => lut_sig <= to_unsigned(integer(my_rom(3176)),16);
when x"c69" => lut_sig <= to_unsigned(integer(my_rom(3177)),16);
when x"c6a" => lut_sig <= to_unsigned(integer(my_rom(3178)),16);
when x"c6b" => lut_sig <= to_unsigned(integer(my_rom(3179)),16);
when x"c6c" => lut_sig <= to_unsigned(integer(my_rom(3180)),16);
when x"c6d" => lut_sig <= to_unsigned(integer(my_rom(3181)),16);
when x"c6e" => lut_sig <= to_unsigned(integer(my_rom(3182)),16);
when x"c6f" => lut_sig <= to_unsigned(integer(my_rom(3183)),16);
when x"c70" => lut_sig <= to_unsigned(integer(my_rom(3184)),16);
when x"c71" => lut_sig <= to_unsigned(integer(my_rom(3185)),16);
when x"c72" => lut_sig <= to_unsigned(integer(my_rom(3186)),16);
when x"c73" => lut_sig <= to_unsigned(integer(my_rom(3187)),16);
when x"c74" => lut_sig <= to_unsigned(integer(my_rom(3188)),16);
when x"c75" => lut_sig <= to_unsigned(integer(my_rom(3189)),16);
when x"c76" => lut_sig <= to_unsigned(integer(my_rom(3190)),16);
when x"c77" => lut_sig <= to_unsigned(integer(my_rom(3191)),16);
when x"c78" => lut_sig <= to_unsigned(integer(my_rom(3192)),16);
when x"c79" => lut_sig <= to_unsigned(integer(my_rom(3193)),16);
when x"c7a" => lut_sig <= to_unsigned(integer(my_rom(3194)),16);
when x"c7b" => lut_sig <= to_unsigned(integer(my_rom(3195)),16);
when x"c7c" => lut_sig <= to_unsigned(integer(my_rom(3196)),16);
when x"c7d" => lut_sig <= to_unsigned(integer(my_rom(3197)),16);
when x"c7e" => lut_sig <= to_unsigned(integer(my_rom(3198)),16);
when x"c7f" => lut_sig <= to_unsigned(integer(my_rom(3199)),16);
when x"c80" => lut_sig <= to_unsigned(integer(my_rom(3200)),16);
when x"c81" => lut_sig <= to_unsigned(integer(my_rom(3201)),16);
when x"c82" => lut_sig <= to_unsigned(integer(my_rom(3202)),16);
when x"c83" => lut_sig <= to_unsigned(integer(my_rom(3203)),16);
when x"c84" => lut_sig <= to_unsigned(integer(my_rom(3204)),16);
when x"c85" => lut_sig <= to_unsigned(integer(my_rom(3205)),16);
when x"c86" => lut_sig <= to_unsigned(integer(my_rom(3206)),16);
when x"c87" => lut_sig <= to_unsigned(integer(my_rom(3207)),16);
when x"c88" => lut_sig <= to_unsigned(integer(my_rom(3208)),16);
when x"c89" => lut_sig <= to_unsigned(integer(my_rom(3209)),16);
when x"c8a" => lut_sig <= to_unsigned(integer(my_rom(3210)),16);
when x"c8b" => lut_sig <= to_unsigned(integer(my_rom(3211)),16);
when x"c8c" => lut_sig <= to_unsigned(integer(my_rom(3212)),16);
when x"c8d" => lut_sig <= to_unsigned(integer(my_rom(3213)),16);
when x"c8e" => lut_sig <= to_unsigned(integer(my_rom(3214)),16);
when x"c8f" => lut_sig <= to_unsigned(integer(my_rom(3215)),16);
when x"c90" => lut_sig <= to_unsigned(integer(my_rom(3216)),16);
when x"c91" => lut_sig <= to_unsigned(integer(my_rom(3217)),16);
when x"c92" => lut_sig <= to_unsigned(integer(my_rom(3218)),16);
when x"c93" => lut_sig <= to_unsigned(integer(my_rom(3219)),16);
when x"c94" => lut_sig <= to_unsigned(integer(my_rom(3220)),16);
when x"c95" => lut_sig <= to_unsigned(integer(my_rom(3221)),16);
when x"c96" => lut_sig <= to_unsigned(integer(my_rom(3222)),16);
when x"c97" => lut_sig <= to_unsigned(integer(my_rom(3223)),16);
when x"c98" => lut_sig <= to_unsigned(integer(my_rom(3224)),16);
when x"c99" => lut_sig <= to_unsigned(integer(my_rom(3225)),16);
when x"c9a" => lut_sig <= to_unsigned(integer(my_rom(3226)),16);
when x"c9b" => lut_sig <= to_unsigned(integer(my_rom(3227)),16);
when x"c9c" => lut_sig <= to_unsigned(integer(my_rom(3228)),16);
when x"c9d" => lut_sig <= to_unsigned(integer(my_rom(3229)),16);
when x"c9e" => lut_sig <= to_unsigned(integer(my_rom(3230)),16);
when x"c9f" => lut_sig <= to_unsigned(integer(my_rom(3231)),16);
when x"ca0" => lut_sig <= to_unsigned(integer(my_rom(3232)),16);
when x"ca1" => lut_sig <= to_unsigned(integer(my_rom(3233)),16);
when x"ca2" => lut_sig <= to_unsigned(integer(my_rom(3234)),16);
when x"ca3" => lut_sig <= to_unsigned(integer(my_rom(3235)),16);
when x"ca4" => lut_sig <= to_unsigned(integer(my_rom(3236)),16);
when x"ca5" => lut_sig <= to_unsigned(integer(my_rom(3237)),16);
when x"ca6" => lut_sig <= to_unsigned(integer(my_rom(3238)),16);
when x"ca7" => lut_sig <= to_unsigned(integer(my_rom(3239)),16);
when x"ca8" => lut_sig <= to_unsigned(integer(my_rom(3240)),16);
when x"ca9" => lut_sig <= to_unsigned(integer(my_rom(3241)),16);
when x"caa" => lut_sig <= to_unsigned(integer(my_rom(3242)),16);
when x"cab" => lut_sig <= to_unsigned(integer(my_rom(3243)),16);
when x"cac" => lut_sig <= to_unsigned(integer(my_rom(3244)),16);
when x"cad" => lut_sig <= to_unsigned(integer(my_rom(3245)),16);
when x"cae" => lut_sig <= to_unsigned(integer(my_rom(3246)),16);
when x"caf" => lut_sig <= to_unsigned(integer(my_rom(3247)),16);
when x"cb0" => lut_sig <= to_unsigned(integer(my_rom(3248)),16);
when x"cb1" => lut_sig <= to_unsigned(integer(my_rom(3249)),16);
when x"cb2" => lut_sig <= to_unsigned(integer(my_rom(3250)),16);
when x"cb3" => lut_sig <= to_unsigned(integer(my_rom(3251)),16);
when x"cb4" => lut_sig <= to_unsigned(integer(my_rom(3252)),16);
when x"cb5" => lut_sig <= to_unsigned(integer(my_rom(3253)),16);
when x"cb6" => lut_sig <= to_unsigned(integer(my_rom(3254)),16);
when x"cb7" => lut_sig <= to_unsigned(integer(my_rom(3255)),16);
when x"cb8" => lut_sig <= to_unsigned(integer(my_rom(3256)),16);
when x"cb9" => lut_sig <= to_unsigned(integer(my_rom(3257)),16);
when x"cba" => lut_sig <= to_unsigned(integer(my_rom(3258)),16);
when x"cbb" => lut_sig <= to_unsigned(integer(my_rom(3259)),16);
when x"cbc" => lut_sig <= to_unsigned(integer(my_rom(3260)),16);
when x"cbd" => lut_sig <= to_unsigned(integer(my_rom(3261)),16);
when x"cbe" => lut_sig <= to_unsigned(integer(my_rom(3262)),16);
when x"cbf" => lut_sig <= to_unsigned(integer(my_rom(3263)),16);
when x"cc0" => lut_sig <= to_unsigned(integer(my_rom(3264)),16);
when x"cc1" => lut_sig <= to_unsigned(integer(my_rom(3265)),16);
when x"cc2" => lut_sig <= to_unsigned(integer(my_rom(3266)),16);
when x"cc3" => lut_sig <= to_unsigned(integer(my_rom(3267)),16);
when x"cc4" => lut_sig <= to_unsigned(integer(my_rom(3268)),16);
when x"cc5" => lut_sig <= to_unsigned(integer(my_rom(3269)),16);
when x"cc6" => lut_sig <= to_unsigned(integer(my_rom(3270)),16);
when x"cc7" => lut_sig <= to_unsigned(integer(my_rom(3271)),16);
when x"cc8" => lut_sig <= to_unsigned(integer(my_rom(3272)),16);
when x"cc9" => lut_sig <= to_unsigned(integer(my_rom(3273)),16);
when x"cca" => lut_sig <= to_unsigned(integer(my_rom(3274)),16);
when x"ccb" => lut_sig <= to_unsigned(integer(my_rom(3275)),16);
when x"ccc" => lut_sig <= to_unsigned(integer(my_rom(3276)),16);
when x"ccd" => lut_sig <= to_unsigned(integer(my_rom(3277)),16);
when x"cce" => lut_sig <= to_unsigned(integer(my_rom(3278)),16);
when x"ccf" => lut_sig <= to_unsigned(integer(my_rom(3279)),16);
when x"cd0" => lut_sig <= to_unsigned(integer(my_rom(3280)),16);
when x"cd1" => lut_sig <= to_unsigned(integer(my_rom(3281)),16);
when x"cd2" => lut_sig <= to_unsigned(integer(my_rom(3282)),16);
when x"cd3" => lut_sig <= to_unsigned(integer(my_rom(3283)),16);
when x"cd4" => lut_sig <= to_unsigned(integer(my_rom(3284)),16);
when x"cd5" => lut_sig <= to_unsigned(integer(my_rom(3285)),16);
when x"cd6" => lut_sig <= to_unsigned(integer(my_rom(3286)),16);
when x"cd7" => lut_sig <= to_unsigned(integer(my_rom(3287)),16);
when x"cd8" => lut_sig <= to_unsigned(integer(my_rom(3288)),16);
when x"cd9" => lut_sig <= to_unsigned(integer(my_rom(3289)),16);
when x"cda" => lut_sig <= to_unsigned(integer(my_rom(3290)),16);
when x"cdb" => lut_sig <= to_unsigned(integer(my_rom(3291)),16);
when x"cdc" => lut_sig <= to_unsigned(integer(my_rom(3292)),16);
when x"cdd" => lut_sig <= to_unsigned(integer(my_rom(3293)),16);
when x"cde" => lut_sig <= to_unsigned(integer(my_rom(3294)),16);
when x"cdf" => lut_sig <= to_unsigned(integer(my_rom(3295)),16);
when x"ce0" => lut_sig <= to_unsigned(integer(my_rom(3296)),16);
when x"ce1" => lut_sig <= to_unsigned(integer(my_rom(3297)),16);
when x"ce2" => lut_sig <= to_unsigned(integer(my_rom(3298)),16);
when x"ce3" => lut_sig <= to_unsigned(integer(my_rom(3299)),16);
when x"ce4" => lut_sig <= to_unsigned(integer(my_rom(3300)),16);
when x"ce5" => lut_sig <= to_unsigned(integer(my_rom(3301)),16);
when x"ce6" => lut_sig <= to_unsigned(integer(my_rom(3302)),16);
when x"ce7" => lut_sig <= to_unsigned(integer(my_rom(3303)),16);
when x"ce8" => lut_sig <= to_unsigned(integer(my_rom(3304)),16);
when x"ce9" => lut_sig <= to_unsigned(integer(my_rom(3305)),16);
when x"cea" => lut_sig <= to_unsigned(integer(my_rom(3306)),16);
when x"ceb" => lut_sig <= to_unsigned(integer(my_rom(3307)),16);
when x"cec" => lut_sig <= to_unsigned(integer(my_rom(3308)),16);
when x"ced" => lut_sig <= to_unsigned(integer(my_rom(3309)),16);
when x"cee" => lut_sig <= to_unsigned(integer(my_rom(3310)),16);
when x"cef" => lut_sig <= to_unsigned(integer(my_rom(3311)),16);
when x"cf0" => lut_sig <= to_unsigned(integer(my_rom(3312)),16);
when x"cf1" => lut_sig <= to_unsigned(integer(my_rom(3313)),16);
when x"cf2" => lut_sig <= to_unsigned(integer(my_rom(3314)),16);
when x"cf3" => lut_sig <= to_unsigned(integer(my_rom(3315)),16);
when x"cf4" => lut_sig <= to_unsigned(integer(my_rom(3316)),16);
when x"cf5" => lut_sig <= to_unsigned(integer(my_rom(3317)),16);
when x"cf6" => lut_sig <= to_unsigned(integer(my_rom(3318)),16);
when x"cf7" => lut_sig <= to_unsigned(integer(my_rom(3319)),16);
when x"cf8" => lut_sig <= to_unsigned(integer(my_rom(3320)),16);
when x"cf9" => lut_sig <= to_unsigned(integer(my_rom(3321)),16);
when x"cfa" => lut_sig <= to_unsigned(integer(my_rom(3322)),16);
when x"cfb" => lut_sig <= to_unsigned(integer(my_rom(3323)),16);
when x"cfc" => lut_sig <= to_unsigned(integer(my_rom(3324)),16);
when x"cfd" => lut_sig <= to_unsigned(integer(my_rom(3325)),16);
when x"cfe" => lut_sig <= to_unsigned(integer(my_rom(3326)),16);
when x"cff" => lut_sig <= to_unsigned(integer(my_rom(3327)),16);
when x"d00" => lut_sig <= to_unsigned(integer(my_rom(3328)),16);
when x"d01" => lut_sig <= to_unsigned(integer(my_rom(3329)),16);
when x"d02" => lut_sig <= to_unsigned(integer(my_rom(3330)),16);
when x"d03" => lut_sig <= to_unsigned(integer(my_rom(3331)),16);
when x"d04" => lut_sig <= to_unsigned(integer(my_rom(3332)),16);
when x"d05" => lut_sig <= to_unsigned(integer(my_rom(3333)),16);
when x"d06" => lut_sig <= to_unsigned(integer(my_rom(3334)),16);
when x"d07" => lut_sig <= to_unsigned(integer(my_rom(3335)),16);
when x"d08" => lut_sig <= to_unsigned(integer(my_rom(3336)),16);
when x"d09" => lut_sig <= to_unsigned(integer(my_rom(3337)),16);
when x"d0a" => lut_sig <= to_unsigned(integer(my_rom(3338)),16);
when x"d0b" => lut_sig <= to_unsigned(integer(my_rom(3339)),16);
when x"d0c" => lut_sig <= to_unsigned(integer(my_rom(3340)),16);
when x"d0d" => lut_sig <= to_unsigned(integer(my_rom(3341)),16);
when x"d0e" => lut_sig <= to_unsigned(integer(my_rom(3342)),16);
when x"d0f" => lut_sig <= to_unsigned(integer(my_rom(3343)),16);
when x"d10" => lut_sig <= to_unsigned(integer(my_rom(3344)),16);
when x"d11" => lut_sig <= to_unsigned(integer(my_rom(3345)),16);
when x"d12" => lut_sig <= to_unsigned(integer(my_rom(3346)),16);
when x"d13" => lut_sig <= to_unsigned(integer(my_rom(3347)),16);
when x"d14" => lut_sig <= to_unsigned(integer(my_rom(3348)),16);
when x"d15" => lut_sig <= to_unsigned(integer(my_rom(3349)),16);
when x"d16" => lut_sig <= to_unsigned(integer(my_rom(3350)),16);
when x"d17" => lut_sig <= to_unsigned(integer(my_rom(3351)),16);
when x"d18" => lut_sig <= to_unsigned(integer(my_rom(3352)),16);
when x"d19" => lut_sig <= to_unsigned(integer(my_rom(3353)),16);
when x"d1a" => lut_sig <= to_unsigned(integer(my_rom(3354)),16);
when x"d1b" => lut_sig <= to_unsigned(integer(my_rom(3355)),16);
when x"d1c" => lut_sig <= to_unsigned(integer(my_rom(3356)),16);
when x"d1d" => lut_sig <= to_unsigned(integer(my_rom(3357)),16);
when x"d1e" => lut_sig <= to_unsigned(integer(my_rom(3358)),16);
when x"d1f" => lut_sig <= to_unsigned(integer(my_rom(3359)),16);
when x"d20" => lut_sig <= to_unsigned(integer(my_rom(3360)),16);
when x"d21" => lut_sig <= to_unsigned(integer(my_rom(3361)),16);
when x"d22" => lut_sig <= to_unsigned(integer(my_rom(3362)),16);
when x"d23" => lut_sig <= to_unsigned(integer(my_rom(3363)),16);
when x"d24" => lut_sig <= to_unsigned(integer(my_rom(3364)),16);
when x"d25" => lut_sig <= to_unsigned(integer(my_rom(3365)),16);
when x"d26" => lut_sig <= to_unsigned(integer(my_rom(3366)),16);
when x"d27" => lut_sig <= to_unsigned(integer(my_rom(3367)),16);
when x"d28" => lut_sig <= to_unsigned(integer(my_rom(3368)),16);
when x"d29" => lut_sig <= to_unsigned(integer(my_rom(3369)),16);
when x"d2a" => lut_sig <= to_unsigned(integer(my_rom(3370)),16);
when x"d2b" => lut_sig <= to_unsigned(integer(my_rom(3371)),16);
when x"d2c" => lut_sig <= to_unsigned(integer(my_rom(3372)),16);
when x"d2d" => lut_sig <= to_unsigned(integer(my_rom(3373)),16);
when x"d2e" => lut_sig <= to_unsigned(integer(my_rom(3374)),16);
when x"d2f" => lut_sig <= to_unsigned(integer(my_rom(3375)),16);
when x"d30" => lut_sig <= to_unsigned(integer(my_rom(3376)),16);
when x"d31" => lut_sig <= to_unsigned(integer(my_rom(3377)),16);
when x"d32" => lut_sig <= to_unsigned(integer(my_rom(3378)),16);
when x"d33" => lut_sig <= to_unsigned(integer(my_rom(3379)),16);
when x"d34" => lut_sig <= to_unsigned(integer(my_rom(3380)),16);
when x"d35" => lut_sig <= to_unsigned(integer(my_rom(3381)),16);
when x"d36" => lut_sig <= to_unsigned(integer(my_rom(3382)),16);
when x"d37" => lut_sig <= to_unsigned(integer(my_rom(3383)),16);
when x"d38" => lut_sig <= to_unsigned(integer(my_rom(3384)),16);
when x"d39" => lut_sig <= to_unsigned(integer(my_rom(3385)),16);
when x"d3a" => lut_sig <= to_unsigned(integer(my_rom(3386)),16);
when x"d3b" => lut_sig <= to_unsigned(integer(my_rom(3387)),16);
when x"d3c" => lut_sig <= to_unsigned(integer(my_rom(3388)),16);
when x"d3d" => lut_sig <= to_unsigned(integer(my_rom(3389)),16);
when x"d3e" => lut_sig <= to_unsigned(integer(my_rom(3390)),16);
when x"d3f" => lut_sig <= to_unsigned(integer(my_rom(3391)),16);
when x"d40" => lut_sig <= to_unsigned(integer(my_rom(3392)),16);
when x"d41" => lut_sig <= to_unsigned(integer(my_rom(3393)),16);
when x"d42" => lut_sig <= to_unsigned(integer(my_rom(3394)),16);
when x"d43" => lut_sig <= to_unsigned(integer(my_rom(3395)),16);
when x"d44" => lut_sig <= to_unsigned(integer(my_rom(3396)),16);
when x"d45" => lut_sig <= to_unsigned(integer(my_rom(3397)),16);
when x"d46" => lut_sig <= to_unsigned(integer(my_rom(3398)),16);
when x"d47" => lut_sig <= to_unsigned(integer(my_rom(3399)),16);
when x"d48" => lut_sig <= to_unsigned(integer(my_rom(3400)),16);
when x"d49" => lut_sig <= to_unsigned(integer(my_rom(3401)),16);
when x"d4a" => lut_sig <= to_unsigned(integer(my_rom(3402)),16);
when x"d4b" => lut_sig <= to_unsigned(integer(my_rom(3403)),16);
when x"d4c" => lut_sig <= to_unsigned(integer(my_rom(3404)),16);
when x"d4d" => lut_sig <= to_unsigned(integer(my_rom(3405)),16);
when x"d4e" => lut_sig <= to_unsigned(integer(my_rom(3406)),16);
when x"d4f" => lut_sig <= to_unsigned(integer(my_rom(3407)),16);
when x"d50" => lut_sig <= to_unsigned(integer(my_rom(3408)),16);
when x"d51" => lut_sig <= to_unsigned(integer(my_rom(3409)),16);
when x"d52" => lut_sig <= to_unsigned(integer(my_rom(3410)),16);
when x"d53" => lut_sig <= to_unsigned(integer(my_rom(3411)),16);
when x"d54" => lut_sig <= to_unsigned(integer(my_rom(3412)),16);
when x"d55" => lut_sig <= to_unsigned(integer(my_rom(3413)),16);
when x"d56" => lut_sig <= to_unsigned(integer(my_rom(3414)),16);
when x"d57" => lut_sig <= to_unsigned(integer(my_rom(3415)),16);
when x"d58" => lut_sig <= to_unsigned(integer(my_rom(3416)),16);
when x"d59" => lut_sig <= to_unsigned(integer(my_rom(3417)),16);
when x"d5a" => lut_sig <= to_unsigned(integer(my_rom(3418)),16);
when x"d5b" => lut_sig <= to_unsigned(integer(my_rom(3419)),16);
when x"d5c" => lut_sig <= to_unsigned(integer(my_rom(3420)),16);
when x"d5d" => lut_sig <= to_unsigned(integer(my_rom(3421)),16);
when x"d5e" => lut_sig <= to_unsigned(integer(my_rom(3422)),16);
when x"d5f" => lut_sig <= to_unsigned(integer(my_rom(3423)),16);
when x"d60" => lut_sig <= to_unsigned(integer(my_rom(3424)),16);
when x"d61" => lut_sig <= to_unsigned(integer(my_rom(3425)),16);
when x"d62" => lut_sig <= to_unsigned(integer(my_rom(3426)),16);
when x"d63" => lut_sig <= to_unsigned(integer(my_rom(3427)),16);
when x"d64" => lut_sig <= to_unsigned(integer(my_rom(3428)),16);
when x"d65" => lut_sig <= to_unsigned(integer(my_rom(3429)),16);
when x"d66" => lut_sig <= to_unsigned(integer(my_rom(3430)),16);
when x"d67" => lut_sig <= to_unsigned(integer(my_rom(3431)),16);
when x"d68" => lut_sig <= to_unsigned(integer(my_rom(3432)),16);
when x"d69" => lut_sig <= to_unsigned(integer(my_rom(3433)),16);
when x"d6a" => lut_sig <= to_unsigned(integer(my_rom(3434)),16);
when x"d6b" => lut_sig <= to_unsigned(integer(my_rom(3435)),16);
when x"d6c" => lut_sig <= to_unsigned(integer(my_rom(3436)),16);
when x"d6d" => lut_sig <= to_unsigned(integer(my_rom(3437)),16);
when x"d6e" => lut_sig <= to_unsigned(integer(my_rom(3438)),16);
when x"d6f" => lut_sig <= to_unsigned(integer(my_rom(3439)),16);
when x"d70" => lut_sig <= to_unsigned(integer(my_rom(3440)),16);
when x"d71" => lut_sig <= to_unsigned(integer(my_rom(3441)),16);
when x"d72" => lut_sig <= to_unsigned(integer(my_rom(3442)),16);
when x"d73" => lut_sig <= to_unsigned(integer(my_rom(3443)),16);
when x"d74" => lut_sig <= to_unsigned(integer(my_rom(3444)),16);
when x"d75" => lut_sig <= to_unsigned(integer(my_rom(3445)),16);
when x"d76" => lut_sig <= to_unsigned(integer(my_rom(3446)),16);
when x"d77" => lut_sig <= to_unsigned(integer(my_rom(3447)),16);
when x"d78" => lut_sig <= to_unsigned(integer(my_rom(3448)),16);
when x"d79" => lut_sig <= to_unsigned(integer(my_rom(3449)),16);
when x"d7a" => lut_sig <= to_unsigned(integer(my_rom(3450)),16);
when x"d7b" => lut_sig <= to_unsigned(integer(my_rom(3451)),16);
when x"d7c" => lut_sig <= to_unsigned(integer(my_rom(3452)),16);
when x"d7d" => lut_sig <= to_unsigned(integer(my_rom(3453)),16);
when x"d7e" => lut_sig <= to_unsigned(integer(my_rom(3454)),16);
when x"d7f" => lut_sig <= to_unsigned(integer(my_rom(3455)),16);
when x"d80" => lut_sig <= to_unsigned(integer(my_rom(3456)),16);
when x"d81" => lut_sig <= to_unsigned(integer(my_rom(3457)),16);
when x"d82" => lut_sig <= to_unsigned(integer(my_rom(3458)),16);
when x"d83" => lut_sig <= to_unsigned(integer(my_rom(3459)),16);
when x"d84" => lut_sig <= to_unsigned(integer(my_rom(3460)),16);
when x"d85" => lut_sig <= to_unsigned(integer(my_rom(3461)),16);
when x"d86" => lut_sig <= to_unsigned(integer(my_rom(3462)),16);
when x"d87" => lut_sig <= to_unsigned(integer(my_rom(3463)),16);
when x"d88" => lut_sig <= to_unsigned(integer(my_rom(3464)),16);
when x"d89" => lut_sig <= to_unsigned(integer(my_rom(3465)),16);
when x"d8a" => lut_sig <= to_unsigned(integer(my_rom(3466)),16);
when x"d8b" => lut_sig <= to_unsigned(integer(my_rom(3467)),16);
when x"d8c" => lut_sig <= to_unsigned(integer(my_rom(3468)),16);
when x"d8d" => lut_sig <= to_unsigned(integer(my_rom(3469)),16);
when x"d8e" => lut_sig <= to_unsigned(integer(my_rom(3470)),16);
when x"d8f" => lut_sig <= to_unsigned(integer(my_rom(3471)),16);
when x"d90" => lut_sig <= to_unsigned(integer(my_rom(3472)),16);
when x"d91" => lut_sig <= to_unsigned(integer(my_rom(3473)),16);
when x"d92" => lut_sig <= to_unsigned(integer(my_rom(3474)),16);
when x"d93" => lut_sig <= to_unsigned(integer(my_rom(3475)),16);
when x"d94" => lut_sig <= to_unsigned(integer(my_rom(3476)),16);
when x"d95" => lut_sig <= to_unsigned(integer(my_rom(3477)),16);
when x"d96" => lut_sig <= to_unsigned(integer(my_rom(3478)),16);
when x"d97" => lut_sig <= to_unsigned(integer(my_rom(3479)),16);
when x"d98" => lut_sig <= to_unsigned(integer(my_rom(3480)),16);
when x"d99" => lut_sig <= to_unsigned(integer(my_rom(3481)),16);
when x"d9a" => lut_sig <= to_unsigned(integer(my_rom(3482)),16);
when x"d9b" => lut_sig <= to_unsigned(integer(my_rom(3483)),16);
when x"d9c" => lut_sig <= to_unsigned(integer(my_rom(3484)),16);
when x"d9d" => lut_sig <= to_unsigned(integer(my_rom(3485)),16);
when x"d9e" => lut_sig <= to_unsigned(integer(my_rom(3486)),16);
when x"d9f" => lut_sig <= to_unsigned(integer(my_rom(3487)),16);
when x"da0" => lut_sig <= to_unsigned(integer(my_rom(3488)),16);
when x"da1" => lut_sig <= to_unsigned(integer(my_rom(3489)),16);
when x"da2" => lut_sig <= to_unsigned(integer(my_rom(3490)),16);
when x"da3" => lut_sig <= to_unsigned(integer(my_rom(3491)),16);
when x"da4" => lut_sig <= to_unsigned(integer(my_rom(3492)),16);
when x"da5" => lut_sig <= to_unsigned(integer(my_rom(3493)),16);
when x"da6" => lut_sig <= to_unsigned(integer(my_rom(3494)),16);
when x"da7" => lut_sig <= to_unsigned(integer(my_rom(3495)),16);
when x"da8" => lut_sig <= to_unsigned(integer(my_rom(3496)),16);
when x"da9" => lut_sig <= to_unsigned(integer(my_rom(3497)),16);
when x"daa" => lut_sig <= to_unsigned(integer(my_rom(3498)),16);
when x"dab" => lut_sig <= to_unsigned(integer(my_rom(3499)),16);
when x"dac" => lut_sig <= to_unsigned(integer(my_rom(3500)),16);
when x"dad" => lut_sig <= to_unsigned(integer(my_rom(3501)),16);
when x"dae" => lut_sig <= to_unsigned(integer(my_rom(3502)),16);
when x"daf" => lut_sig <= to_unsigned(integer(my_rom(3503)),16);
when x"db0" => lut_sig <= to_unsigned(integer(my_rom(3504)),16);
when x"db1" => lut_sig <= to_unsigned(integer(my_rom(3505)),16);
when x"db2" => lut_sig <= to_unsigned(integer(my_rom(3506)),16);
when x"db3" => lut_sig <= to_unsigned(integer(my_rom(3507)),16);
when x"db4" => lut_sig <= to_unsigned(integer(my_rom(3508)),16);
when x"db5" => lut_sig <= to_unsigned(integer(my_rom(3509)),16);
when x"db6" => lut_sig <= to_unsigned(integer(my_rom(3510)),16);
when x"db7" => lut_sig <= to_unsigned(integer(my_rom(3511)),16);
when x"db8" => lut_sig <= to_unsigned(integer(my_rom(3512)),16);
when x"db9" => lut_sig <= to_unsigned(integer(my_rom(3513)),16);
when x"dba" => lut_sig <= to_unsigned(integer(my_rom(3514)),16);
when x"dbb" => lut_sig <= to_unsigned(integer(my_rom(3515)),16);
when x"dbc" => lut_sig <= to_unsigned(integer(my_rom(3516)),16);
when x"dbd" => lut_sig <= to_unsigned(integer(my_rom(3517)),16);
when x"dbe" => lut_sig <= to_unsigned(integer(my_rom(3518)),16);
when x"dbf" => lut_sig <= to_unsigned(integer(my_rom(3519)),16);
when x"dc0" => lut_sig <= to_unsigned(integer(my_rom(3520)),16);
when x"dc1" => lut_sig <= to_unsigned(integer(my_rom(3521)),16);
when x"dc2" => lut_sig <= to_unsigned(integer(my_rom(3522)),16);
when x"dc3" => lut_sig <= to_unsigned(integer(my_rom(3523)),16);
when x"dc4" => lut_sig <= to_unsigned(integer(my_rom(3524)),16);
when x"dc5" => lut_sig <= to_unsigned(integer(my_rom(3525)),16);
when x"dc6" => lut_sig <= to_unsigned(integer(my_rom(3526)),16);
when x"dc7" => lut_sig <= to_unsigned(integer(my_rom(3527)),16);
when x"dc8" => lut_sig <= to_unsigned(integer(my_rom(3528)),16);
when x"dc9" => lut_sig <= to_unsigned(integer(my_rom(3529)),16);
when x"dca" => lut_sig <= to_unsigned(integer(my_rom(3530)),16);
when x"dcb" => lut_sig <= to_unsigned(integer(my_rom(3531)),16);
when x"dcc" => lut_sig <= to_unsigned(integer(my_rom(3532)),16);
when x"dcd" => lut_sig <= to_unsigned(integer(my_rom(3533)),16);
when x"dce" => lut_sig <= to_unsigned(integer(my_rom(3534)),16);
when x"dcf" => lut_sig <= to_unsigned(integer(my_rom(3535)),16);
when x"dd0" => lut_sig <= to_unsigned(integer(my_rom(3536)),16);
when x"dd1" => lut_sig <= to_unsigned(integer(my_rom(3537)),16);
when x"dd2" => lut_sig <= to_unsigned(integer(my_rom(3538)),16);
when x"dd3" => lut_sig <= to_unsigned(integer(my_rom(3539)),16);
when x"dd4" => lut_sig <= to_unsigned(integer(my_rom(3540)),16);
when x"dd5" => lut_sig <= to_unsigned(integer(my_rom(3541)),16);
when x"dd6" => lut_sig <= to_unsigned(integer(my_rom(3542)),16);
when x"dd7" => lut_sig <= to_unsigned(integer(my_rom(3543)),16);
when x"dd8" => lut_sig <= to_unsigned(integer(my_rom(3544)),16);
when x"dd9" => lut_sig <= to_unsigned(integer(my_rom(3545)),16);
when x"dda" => lut_sig <= to_unsigned(integer(my_rom(3546)),16);
when x"ddb" => lut_sig <= to_unsigned(integer(my_rom(3547)),16);
when x"ddc" => lut_sig <= to_unsigned(integer(my_rom(3548)),16);
when x"ddd" => lut_sig <= to_unsigned(integer(my_rom(3549)),16);
when x"dde" => lut_sig <= to_unsigned(integer(my_rom(3550)),16);
when x"ddf" => lut_sig <= to_unsigned(integer(my_rom(3551)),16);
when x"de0" => lut_sig <= to_unsigned(integer(my_rom(3552)),16);
when x"de1" => lut_sig <= to_unsigned(integer(my_rom(3553)),16);
when x"de2" => lut_sig <= to_unsigned(integer(my_rom(3554)),16);
when x"de3" => lut_sig <= to_unsigned(integer(my_rom(3555)),16);
when x"de4" => lut_sig <= to_unsigned(integer(my_rom(3556)),16);
when x"de5" => lut_sig <= to_unsigned(integer(my_rom(3557)),16);
when x"de6" => lut_sig <= to_unsigned(integer(my_rom(3558)),16);
when x"de7" => lut_sig <= to_unsigned(integer(my_rom(3559)),16);
when x"de8" => lut_sig <= to_unsigned(integer(my_rom(3560)),16);
when x"de9" => lut_sig <= to_unsigned(integer(my_rom(3561)),16);
when x"dea" => lut_sig <= to_unsigned(integer(my_rom(3562)),16);
when x"deb" => lut_sig <= to_unsigned(integer(my_rom(3563)),16);
when x"dec" => lut_sig <= to_unsigned(integer(my_rom(3564)),16);
when x"ded" => lut_sig <= to_unsigned(integer(my_rom(3565)),16);
when x"dee" => lut_sig <= to_unsigned(integer(my_rom(3566)),16);
when x"def" => lut_sig <= to_unsigned(integer(my_rom(3567)),16);
when x"df0" => lut_sig <= to_unsigned(integer(my_rom(3568)),16);
when x"df1" => lut_sig <= to_unsigned(integer(my_rom(3569)),16);
when x"df2" => lut_sig <= to_unsigned(integer(my_rom(3570)),16);
when x"df3" => lut_sig <= to_unsigned(integer(my_rom(3571)),16);
when x"df4" => lut_sig <= to_unsigned(integer(my_rom(3572)),16);
when x"df5" => lut_sig <= to_unsigned(integer(my_rom(3573)),16);
when x"df6" => lut_sig <= to_unsigned(integer(my_rom(3574)),16);
when x"df7" => lut_sig <= to_unsigned(integer(my_rom(3575)),16);
when x"df8" => lut_sig <= to_unsigned(integer(my_rom(3576)),16);
when x"df9" => lut_sig <= to_unsigned(integer(my_rom(3577)),16);
when x"dfa" => lut_sig <= to_unsigned(integer(my_rom(3578)),16);
when x"dfb" => lut_sig <= to_unsigned(integer(my_rom(3579)),16);
when x"dfc" => lut_sig <= to_unsigned(integer(my_rom(3580)),16);
when x"dfd" => lut_sig <= to_unsigned(integer(my_rom(3581)),16);
when x"dfe" => lut_sig <= to_unsigned(integer(my_rom(3582)),16);
when x"dff" => lut_sig <= to_unsigned(integer(my_rom(3583)),16);
when x"e00" => lut_sig <= to_unsigned(integer(my_rom(3584)),16);
when x"e01" => lut_sig <= to_unsigned(integer(my_rom(3585)),16);
when x"e02" => lut_sig <= to_unsigned(integer(my_rom(3586)),16);
when x"e03" => lut_sig <= to_unsigned(integer(my_rom(3587)),16);
when x"e04" => lut_sig <= to_unsigned(integer(my_rom(3588)),16);
when x"e05" => lut_sig <= to_unsigned(integer(my_rom(3589)),16);
when x"e06" => lut_sig <= to_unsigned(integer(my_rom(3590)),16);
when x"e07" => lut_sig <= to_unsigned(integer(my_rom(3591)),16);
when x"e08" => lut_sig <= to_unsigned(integer(my_rom(3592)),16);
when x"e09" => lut_sig <= to_unsigned(integer(my_rom(3593)),16);
when x"e0a" => lut_sig <= to_unsigned(integer(my_rom(3594)),16);
when x"e0b" => lut_sig <= to_unsigned(integer(my_rom(3595)),16);
when x"e0c" => lut_sig <= to_unsigned(integer(my_rom(3596)),16);
when x"e0d" => lut_sig <= to_unsigned(integer(my_rom(3597)),16);
when x"e0e" => lut_sig <= to_unsigned(integer(my_rom(3598)),16);
when x"e0f" => lut_sig <= to_unsigned(integer(my_rom(3599)),16);
when x"e10" => lut_sig <= to_unsigned(integer(my_rom(3600)),16);
when x"e11" => lut_sig <= to_unsigned(integer(my_rom(3601)),16);
when x"e12" => lut_sig <= to_unsigned(integer(my_rom(3602)),16);
when x"e13" => lut_sig <= to_unsigned(integer(my_rom(3603)),16);
when x"e14" => lut_sig <= to_unsigned(integer(my_rom(3604)),16);
when x"e15" => lut_sig <= to_unsigned(integer(my_rom(3605)),16);
when x"e16" => lut_sig <= to_unsigned(integer(my_rom(3606)),16);
when x"e17" => lut_sig <= to_unsigned(integer(my_rom(3607)),16);
when x"e18" => lut_sig <= to_unsigned(integer(my_rom(3608)),16);
when x"e19" => lut_sig <= to_unsigned(integer(my_rom(3609)),16);
when x"e1a" => lut_sig <= to_unsigned(integer(my_rom(3610)),16);
when x"e1b" => lut_sig <= to_unsigned(integer(my_rom(3611)),16);
when x"e1c" => lut_sig <= to_unsigned(integer(my_rom(3612)),16);
when x"e1d" => lut_sig <= to_unsigned(integer(my_rom(3613)),16);
when x"e1e" => lut_sig <= to_unsigned(integer(my_rom(3614)),16);
when x"e1f" => lut_sig <= to_unsigned(integer(my_rom(3615)),16);
when x"e20" => lut_sig <= to_unsigned(integer(my_rom(3616)),16);
when x"e21" => lut_sig <= to_unsigned(integer(my_rom(3617)),16);
when x"e22" => lut_sig <= to_unsigned(integer(my_rom(3618)),16);
when x"e23" => lut_sig <= to_unsigned(integer(my_rom(3619)),16);
when x"e24" => lut_sig <= to_unsigned(integer(my_rom(3620)),16);
when x"e25" => lut_sig <= to_unsigned(integer(my_rom(3621)),16);
when x"e26" => lut_sig <= to_unsigned(integer(my_rom(3622)),16);
when x"e27" => lut_sig <= to_unsigned(integer(my_rom(3623)),16);
when x"e28" => lut_sig <= to_unsigned(integer(my_rom(3624)),16);
when x"e29" => lut_sig <= to_unsigned(integer(my_rom(3625)),16);
when x"e2a" => lut_sig <= to_unsigned(integer(my_rom(3626)),16);
when x"e2b" => lut_sig <= to_unsigned(integer(my_rom(3627)),16);
when x"e2c" => lut_sig <= to_unsigned(integer(my_rom(3628)),16);
when x"e2d" => lut_sig <= to_unsigned(integer(my_rom(3629)),16);
when x"e2e" => lut_sig <= to_unsigned(integer(my_rom(3630)),16);
when x"e2f" => lut_sig <= to_unsigned(integer(my_rom(3631)),16);
when x"e30" => lut_sig <= to_unsigned(integer(my_rom(3632)),16);
when x"e31" => lut_sig <= to_unsigned(integer(my_rom(3633)),16);
when x"e32" => lut_sig <= to_unsigned(integer(my_rom(3634)),16);
when x"e33" => lut_sig <= to_unsigned(integer(my_rom(3635)),16);
when x"e34" => lut_sig <= to_unsigned(integer(my_rom(3636)),16);
when x"e35" => lut_sig <= to_unsigned(integer(my_rom(3637)),16);
when x"e36" => lut_sig <= to_unsigned(integer(my_rom(3638)),16);
when x"e37" => lut_sig <= to_unsigned(integer(my_rom(3639)),16);
when x"e38" => lut_sig <= to_unsigned(integer(my_rom(3640)),16);
when x"e39" => lut_sig <= to_unsigned(integer(my_rom(3641)),16);
when x"e3a" => lut_sig <= to_unsigned(integer(my_rom(3642)),16);
when x"e3b" => lut_sig <= to_unsigned(integer(my_rom(3643)),16);
when x"e3c" => lut_sig <= to_unsigned(integer(my_rom(3644)),16);
when x"e3d" => lut_sig <= to_unsigned(integer(my_rom(3645)),16);
when x"e3e" => lut_sig <= to_unsigned(integer(my_rom(3646)),16);
when x"e3f" => lut_sig <= to_unsigned(integer(my_rom(3647)),16);
when x"e40" => lut_sig <= to_unsigned(integer(my_rom(3648)),16);
when x"e41" => lut_sig <= to_unsigned(integer(my_rom(3649)),16);
when x"e42" => lut_sig <= to_unsigned(integer(my_rom(3650)),16);
when x"e43" => lut_sig <= to_unsigned(integer(my_rom(3651)),16);
when x"e44" => lut_sig <= to_unsigned(integer(my_rom(3652)),16);
when x"e45" => lut_sig <= to_unsigned(integer(my_rom(3653)),16);
when x"e46" => lut_sig <= to_unsigned(integer(my_rom(3654)),16);
when x"e47" => lut_sig <= to_unsigned(integer(my_rom(3655)),16);
when x"e48" => lut_sig <= to_unsigned(integer(my_rom(3656)),16);
when x"e49" => lut_sig <= to_unsigned(integer(my_rom(3657)),16);
when x"e4a" => lut_sig <= to_unsigned(integer(my_rom(3658)),16);
when x"e4b" => lut_sig <= to_unsigned(integer(my_rom(3659)),16);
when x"e4c" => lut_sig <= to_unsigned(integer(my_rom(3660)),16);
when x"e4d" => lut_sig <= to_unsigned(integer(my_rom(3661)),16);
when x"e4e" => lut_sig <= to_unsigned(integer(my_rom(3662)),16);
when x"e4f" => lut_sig <= to_unsigned(integer(my_rom(3663)),16);
when x"e50" => lut_sig <= to_unsigned(integer(my_rom(3664)),16);
when x"e51" => lut_sig <= to_unsigned(integer(my_rom(3665)),16);
when x"e52" => lut_sig <= to_unsigned(integer(my_rom(3666)),16);
when x"e53" => lut_sig <= to_unsigned(integer(my_rom(3667)),16);
when x"e54" => lut_sig <= to_unsigned(integer(my_rom(3668)),16);
when x"e55" => lut_sig <= to_unsigned(integer(my_rom(3669)),16);
when x"e56" => lut_sig <= to_unsigned(integer(my_rom(3670)),16);
when x"e57" => lut_sig <= to_unsigned(integer(my_rom(3671)),16);
when x"e58" => lut_sig <= to_unsigned(integer(my_rom(3672)),16);
when x"e59" => lut_sig <= to_unsigned(integer(my_rom(3673)),16);
when x"e5a" => lut_sig <= to_unsigned(integer(my_rom(3674)),16);
when x"e5b" => lut_sig <= to_unsigned(integer(my_rom(3675)),16);
when x"e5c" => lut_sig <= to_unsigned(integer(my_rom(3676)),16);
when x"e5d" => lut_sig <= to_unsigned(integer(my_rom(3677)),16);
when x"e5e" => lut_sig <= to_unsigned(integer(my_rom(3678)),16);
when x"e5f" => lut_sig <= to_unsigned(integer(my_rom(3679)),16);
when x"e60" => lut_sig <= to_unsigned(integer(my_rom(3680)),16);
when x"e61" => lut_sig <= to_unsigned(integer(my_rom(3681)),16);
when x"e62" => lut_sig <= to_unsigned(integer(my_rom(3682)),16);
when x"e63" => lut_sig <= to_unsigned(integer(my_rom(3683)),16);
when x"e64" => lut_sig <= to_unsigned(integer(my_rom(3684)),16);
when x"e65" => lut_sig <= to_unsigned(integer(my_rom(3685)),16);
when x"e66" => lut_sig <= to_unsigned(integer(my_rom(3686)),16);
when x"e67" => lut_sig <= to_unsigned(integer(my_rom(3687)),16);
when x"e68" => lut_sig <= to_unsigned(integer(my_rom(3688)),16);
when x"e69" => lut_sig <= to_unsigned(integer(my_rom(3689)),16);
when x"e6a" => lut_sig <= to_unsigned(integer(my_rom(3690)),16);
when x"e6b" => lut_sig <= to_unsigned(integer(my_rom(3691)),16);
when x"e6c" => lut_sig <= to_unsigned(integer(my_rom(3692)),16);
when x"e6d" => lut_sig <= to_unsigned(integer(my_rom(3693)),16);
when x"e6e" => lut_sig <= to_unsigned(integer(my_rom(3694)),16);
when x"e6f" => lut_sig <= to_unsigned(integer(my_rom(3695)),16);
when x"e70" => lut_sig <= to_unsigned(integer(my_rom(3696)),16);
when x"e71" => lut_sig <= to_unsigned(integer(my_rom(3697)),16);
when x"e72" => lut_sig <= to_unsigned(integer(my_rom(3698)),16);
when x"e73" => lut_sig <= to_unsigned(integer(my_rom(3699)),16);
when x"e74" => lut_sig <= to_unsigned(integer(my_rom(3700)),16);
when x"e75" => lut_sig <= to_unsigned(integer(my_rom(3701)),16);
when x"e76" => lut_sig <= to_unsigned(integer(my_rom(3702)),16);
when x"e77" => lut_sig <= to_unsigned(integer(my_rom(3703)),16);
when x"e78" => lut_sig <= to_unsigned(integer(my_rom(3704)),16);
when x"e79" => lut_sig <= to_unsigned(integer(my_rom(3705)),16);
when x"e7a" => lut_sig <= to_unsigned(integer(my_rom(3706)),16);
when x"e7b" => lut_sig <= to_unsigned(integer(my_rom(3707)),16);
when x"e7c" => lut_sig <= to_unsigned(integer(my_rom(3708)),16);
when x"e7d" => lut_sig <= to_unsigned(integer(my_rom(3709)),16);
when x"e7e" => lut_sig <= to_unsigned(integer(my_rom(3710)),16);
when x"e7f" => lut_sig <= to_unsigned(integer(my_rom(3711)),16);
when x"e80" => lut_sig <= to_unsigned(integer(my_rom(3712)),16);
when x"e81" => lut_sig <= to_unsigned(integer(my_rom(3713)),16);
when x"e82" => lut_sig <= to_unsigned(integer(my_rom(3714)),16);
when x"e83" => lut_sig <= to_unsigned(integer(my_rom(3715)),16);
when x"e84" => lut_sig <= to_unsigned(integer(my_rom(3716)),16);
when x"e85" => lut_sig <= to_unsigned(integer(my_rom(3717)),16);
when x"e86" => lut_sig <= to_unsigned(integer(my_rom(3718)),16);
when x"e87" => lut_sig <= to_unsigned(integer(my_rom(3719)),16);
when x"e88" => lut_sig <= to_unsigned(integer(my_rom(3720)),16);
when x"e89" => lut_sig <= to_unsigned(integer(my_rom(3721)),16);
when x"e8a" => lut_sig <= to_unsigned(integer(my_rom(3722)),16);
when x"e8b" => lut_sig <= to_unsigned(integer(my_rom(3723)),16);
when x"e8c" => lut_sig <= to_unsigned(integer(my_rom(3724)),16);
when x"e8d" => lut_sig <= to_unsigned(integer(my_rom(3725)),16);
when x"e8e" => lut_sig <= to_unsigned(integer(my_rom(3726)),16);
when x"e8f" => lut_sig <= to_unsigned(integer(my_rom(3727)),16);
when x"e90" => lut_sig <= to_unsigned(integer(my_rom(3728)),16);
when x"e91" => lut_sig <= to_unsigned(integer(my_rom(3729)),16);
when x"e92" => lut_sig <= to_unsigned(integer(my_rom(3730)),16);
when x"e93" => lut_sig <= to_unsigned(integer(my_rom(3731)),16);
when x"e94" => lut_sig <= to_unsigned(integer(my_rom(3732)),16);
when x"e95" => lut_sig <= to_unsigned(integer(my_rom(3733)),16);
when x"e96" => lut_sig <= to_unsigned(integer(my_rom(3734)),16);
when x"e97" => lut_sig <= to_unsigned(integer(my_rom(3735)),16);
when x"e98" => lut_sig <= to_unsigned(integer(my_rom(3736)),16);
when x"e99" => lut_sig <= to_unsigned(integer(my_rom(3737)),16);
when x"e9a" => lut_sig <= to_unsigned(integer(my_rom(3738)),16);
when x"e9b" => lut_sig <= to_unsigned(integer(my_rom(3739)),16);
when x"e9c" => lut_sig <= to_unsigned(integer(my_rom(3740)),16);
when x"e9d" => lut_sig <= to_unsigned(integer(my_rom(3741)),16);
when x"e9e" => lut_sig <= to_unsigned(integer(my_rom(3742)),16);
when x"e9f" => lut_sig <= to_unsigned(integer(my_rom(3743)),16);
when x"ea0" => lut_sig <= to_unsigned(integer(my_rom(3744)),16);
when x"ea1" => lut_sig <= to_unsigned(integer(my_rom(3745)),16);
when x"ea2" => lut_sig <= to_unsigned(integer(my_rom(3746)),16);
when x"ea3" => lut_sig <= to_unsigned(integer(my_rom(3747)),16);
when x"ea4" => lut_sig <= to_unsigned(integer(my_rom(3748)),16);
when x"ea5" => lut_sig <= to_unsigned(integer(my_rom(3749)),16);
when x"ea6" => lut_sig <= to_unsigned(integer(my_rom(3750)),16);
when x"ea7" => lut_sig <= to_unsigned(integer(my_rom(3751)),16);
when x"ea8" => lut_sig <= to_unsigned(integer(my_rom(3752)),16);
when x"ea9" => lut_sig <= to_unsigned(integer(my_rom(3753)),16);
when x"eaa" => lut_sig <= to_unsigned(integer(my_rom(3754)),16);
when x"eab" => lut_sig <= to_unsigned(integer(my_rom(3755)),16);
when x"eac" => lut_sig <= to_unsigned(integer(my_rom(3756)),16);
when x"ead" => lut_sig <= to_unsigned(integer(my_rom(3757)),16);
when x"eae" => lut_sig <= to_unsigned(integer(my_rom(3758)),16);
when x"eaf" => lut_sig <= to_unsigned(integer(my_rom(3759)),16);
when x"eb0" => lut_sig <= to_unsigned(integer(my_rom(3760)),16);
when x"eb1" => lut_sig <= to_unsigned(integer(my_rom(3761)),16);
when x"eb2" => lut_sig <= to_unsigned(integer(my_rom(3762)),16);
when x"eb3" => lut_sig <= to_unsigned(integer(my_rom(3763)),16);
when x"eb4" => lut_sig <= to_unsigned(integer(my_rom(3764)),16);
when x"eb5" => lut_sig <= to_unsigned(integer(my_rom(3765)),16);
when x"eb6" => lut_sig <= to_unsigned(integer(my_rom(3766)),16);
when x"eb7" => lut_sig <= to_unsigned(integer(my_rom(3767)),16);
when x"eb8" => lut_sig <= to_unsigned(integer(my_rom(3768)),16);
when x"eb9" => lut_sig <= to_unsigned(integer(my_rom(3769)),16);
when x"eba" => lut_sig <= to_unsigned(integer(my_rom(3770)),16);
when x"ebb" => lut_sig <= to_unsigned(integer(my_rom(3771)),16);
when x"ebc" => lut_sig <= to_unsigned(integer(my_rom(3772)),16);
when x"ebd" => lut_sig <= to_unsigned(integer(my_rom(3773)),16);
when x"ebe" => lut_sig <= to_unsigned(integer(my_rom(3774)),16);
when x"ebf" => lut_sig <= to_unsigned(integer(my_rom(3775)),16);
when x"ec0" => lut_sig <= to_unsigned(integer(my_rom(3776)),16);
when x"ec1" => lut_sig <= to_unsigned(integer(my_rom(3777)),16);
when x"ec2" => lut_sig <= to_unsigned(integer(my_rom(3778)),16);
when x"ec3" => lut_sig <= to_unsigned(integer(my_rom(3779)),16);
when x"ec4" => lut_sig <= to_unsigned(integer(my_rom(3780)),16);
when x"ec5" => lut_sig <= to_unsigned(integer(my_rom(3781)),16);
when x"ec6" => lut_sig <= to_unsigned(integer(my_rom(3782)),16);
when x"ec7" => lut_sig <= to_unsigned(integer(my_rom(3783)),16);
when x"ec8" => lut_sig <= to_unsigned(integer(my_rom(3784)),16);
when x"ec9" => lut_sig <= to_unsigned(integer(my_rom(3785)),16);
when x"eca" => lut_sig <= to_unsigned(integer(my_rom(3786)),16);
when x"ecb" => lut_sig <= to_unsigned(integer(my_rom(3787)),16);
when x"ecc" => lut_sig <= to_unsigned(integer(my_rom(3788)),16);
when x"ecd" => lut_sig <= to_unsigned(integer(my_rom(3789)),16);
when x"ece" => lut_sig <= to_unsigned(integer(my_rom(3790)),16);
when x"ecf" => lut_sig <= to_unsigned(integer(my_rom(3791)),16);
when x"ed0" => lut_sig <= to_unsigned(integer(my_rom(3792)),16);
when x"ed1" => lut_sig <= to_unsigned(integer(my_rom(3793)),16);
when x"ed2" => lut_sig <= to_unsigned(integer(my_rom(3794)),16);
when x"ed3" => lut_sig <= to_unsigned(integer(my_rom(3795)),16);
when x"ed4" => lut_sig <= to_unsigned(integer(my_rom(3796)),16);
when x"ed5" => lut_sig <= to_unsigned(integer(my_rom(3797)),16);
when x"ed6" => lut_sig <= to_unsigned(integer(my_rom(3798)),16);
when x"ed7" => lut_sig <= to_unsigned(integer(my_rom(3799)),16);
when x"ed8" => lut_sig <= to_unsigned(integer(my_rom(3800)),16);
when x"ed9" => lut_sig <= to_unsigned(integer(my_rom(3801)),16);
when x"eda" => lut_sig <= to_unsigned(integer(my_rom(3802)),16);
when x"edb" => lut_sig <= to_unsigned(integer(my_rom(3803)),16);
when x"edc" => lut_sig <= to_unsigned(integer(my_rom(3804)),16);
when x"edd" => lut_sig <= to_unsigned(integer(my_rom(3805)),16);
when x"ede" => lut_sig <= to_unsigned(integer(my_rom(3806)),16);
when x"edf" => lut_sig <= to_unsigned(integer(my_rom(3807)),16);
when x"ee0" => lut_sig <= to_unsigned(integer(my_rom(3808)),16);
when x"ee1" => lut_sig <= to_unsigned(integer(my_rom(3809)),16);
when x"ee2" => lut_sig <= to_unsigned(integer(my_rom(3810)),16);
when x"ee3" => lut_sig <= to_unsigned(integer(my_rom(3811)),16);
when x"ee4" => lut_sig <= to_unsigned(integer(my_rom(3812)),16);
when x"ee5" => lut_sig <= to_unsigned(integer(my_rom(3813)),16);
when x"ee6" => lut_sig <= to_unsigned(integer(my_rom(3814)),16);
when x"ee7" => lut_sig <= to_unsigned(integer(my_rom(3815)),16);
when x"ee8" => lut_sig <= to_unsigned(integer(my_rom(3816)),16);
when x"ee9" => lut_sig <= to_unsigned(integer(my_rom(3817)),16);
when x"eea" => lut_sig <= to_unsigned(integer(my_rom(3818)),16);
when x"eeb" => lut_sig <= to_unsigned(integer(my_rom(3819)),16);
when x"eec" => lut_sig <= to_unsigned(integer(my_rom(3820)),16);
when x"eed" => lut_sig <= to_unsigned(integer(my_rom(3821)),16);
when x"eee" => lut_sig <= to_unsigned(integer(my_rom(3822)),16);
when x"eef" => lut_sig <= to_unsigned(integer(my_rom(3823)),16);
when x"ef0" => lut_sig <= to_unsigned(integer(my_rom(3824)),16);
when x"ef1" => lut_sig <= to_unsigned(integer(my_rom(3825)),16);
when x"ef2" => lut_sig <= to_unsigned(integer(my_rom(3826)),16);
when x"ef3" => lut_sig <= to_unsigned(integer(my_rom(3827)),16);
when x"ef4" => lut_sig <= to_unsigned(integer(my_rom(3828)),16);
when x"ef5" => lut_sig <= to_unsigned(integer(my_rom(3829)),16);
when x"ef6" => lut_sig <= to_unsigned(integer(my_rom(3830)),16);
when x"ef7" => lut_sig <= to_unsigned(integer(my_rom(3831)),16);
when x"ef8" => lut_sig <= to_unsigned(integer(my_rom(3832)),16);
when x"ef9" => lut_sig <= to_unsigned(integer(my_rom(3833)),16);
when x"efa" => lut_sig <= to_unsigned(integer(my_rom(3834)),16);
when x"efb" => lut_sig <= to_unsigned(integer(my_rom(3835)),16);
when x"efc" => lut_sig <= to_unsigned(integer(my_rom(3836)),16);
when x"efd" => lut_sig <= to_unsigned(integer(my_rom(3837)),16);
when x"efe" => lut_sig <= to_unsigned(integer(my_rom(3838)),16);
when x"eff" => lut_sig <= to_unsigned(integer(my_rom(3839)),16);
when x"f00" => lut_sig <= to_unsigned(integer(my_rom(3840)),16);
when x"f01" => lut_sig <= to_unsigned(integer(my_rom(3841)),16);
when x"f02" => lut_sig <= to_unsigned(integer(my_rom(3842)),16);
when x"f03" => lut_sig <= to_unsigned(integer(my_rom(3843)),16);
when x"f04" => lut_sig <= to_unsigned(integer(my_rom(3844)),16);
when x"f05" => lut_sig <= to_unsigned(integer(my_rom(3845)),16);
when x"f06" => lut_sig <= to_unsigned(integer(my_rom(3846)),16);
when x"f07" => lut_sig <= to_unsigned(integer(my_rom(3847)),16);
when x"f08" => lut_sig <= to_unsigned(integer(my_rom(3848)),16);
when x"f09" => lut_sig <= to_unsigned(integer(my_rom(3849)),16);
when x"f0a" => lut_sig <= to_unsigned(integer(my_rom(3850)),16);
when x"f0b" => lut_sig <= to_unsigned(integer(my_rom(3851)),16);
when x"f0c" => lut_sig <= to_unsigned(integer(my_rom(3852)),16);
when x"f0d" => lut_sig <= to_unsigned(integer(my_rom(3853)),16);
when x"f0e" => lut_sig <= to_unsigned(integer(my_rom(3854)),16);
when x"f0f" => lut_sig <= to_unsigned(integer(my_rom(3855)),16);
when x"f10" => lut_sig <= to_unsigned(integer(my_rom(3856)),16);
when x"f11" => lut_sig <= to_unsigned(integer(my_rom(3857)),16);
when x"f12" => lut_sig <= to_unsigned(integer(my_rom(3858)),16);
when x"f13" => lut_sig <= to_unsigned(integer(my_rom(3859)),16);
when x"f14" => lut_sig <= to_unsigned(integer(my_rom(3860)),16);
when x"f15" => lut_sig <= to_unsigned(integer(my_rom(3861)),16);
when x"f16" => lut_sig <= to_unsigned(integer(my_rom(3862)),16);
when x"f17" => lut_sig <= to_unsigned(integer(my_rom(3863)),16);
when x"f18" => lut_sig <= to_unsigned(integer(my_rom(3864)),16);
when x"f19" => lut_sig <= to_unsigned(integer(my_rom(3865)),16);
when x"f1a" => lut_sig <= to_unsigned(integer(my_rom(3866)),16);
when x"f1b" => lut_sig <= to_unsigned(integer(my_rom(3867)),16);
when x"f1c" => lut_sig <= to_unsigned(integer(my_rom(3868)),16);
when x"f1d" => lut_sig <= to_unsigned(integer(my_rom(3869)),16);
when x"f1e" => lut_sig <= to_unsigned(integer(my_rom(3870)),16);
when x"f1f" => lut_sig <= to_unsigned(integer(my_rom(3871)),16);
when x"f20" => lut_sig <= to_unsigned(integer(my_rom(3872)),16);
when x"f21" => lut_sig <= to_unsigned(integer(my_rom(3873)),16);
when x"f22" => lut_sig <= to_unsigned(integer(my_rom(3874)),16);
when x"f23" => lut_sig <= to_unsigned(integer(my_rom(3875)),16);
when x"f24" => lut_sig <= to_unsigned(integer(my_rom(3876)),16);
when x"f25" => lut_sig <= to_unsigned(integer(my_rom(3877)),16);
when x"f26" => lut_sig <= to_unsigned(integer(my_rom(3878)),16);
when x"f27" => lut_sig <= to_unsigned(integer(my_rom(3879)),16);
when x"f28" => lut_sig <= to_unsigned(integer(my_rom(3880)),16);
when x"f29" => lut_sig <= to_unsigned(integer(my_rom(3881)),16);
when x"f2a" => lut_sig <= to_unsigned(integer(my_rom(3882)),16);
when x"f2b" => lut_sig <= to_unsigned(integer(my_rom(3883)),16);
when x"f2c" => lut_sig <= to_unsigned(integer(my_rom(3884)),16);
when x"f2d" => lut_sig <= to_unsigned(integer(my_rom(3885)),16);
when x"f2e" => lut_sig <= to_unsigned(integer(my_rom(3886)),16);
when x"f2f" => lut_sig <= to_unsigned(integer(my_rom(3887)),16);
when x"f30" => lut_sig <= to_unsigned(integer(my_rom(3888)),16);
when x"f31" => lut_sig <= to_unsigned(integer(my_rom(3889)),16);
when x"f32" => lut_sig <= to_unsigned(integer(my_rom(3890)),16);
when x"f33" => lut_sig <= to_unsigned(integer(my_rom(3891)),16);
when x"f34" => lut_sig <= to_unsigned(integer(my_rom(3892)),16);
when x"f35" => lut_sig <= to_unsigned(integer(my_rom(3893)),16);
when x"f36" => lut_sig <= to_unsigned(integer(my_rom(3894)),16);
when x"f37" => lut_sig <= to_unsigned(integer(my_rom(3895)),16);
when x"f38" => lut_sig <= to_unsigned(integer(my_rom(3896)),16);
when x"f39" => lut_sig <= to_unsigned(integer(my_rom(3897)),16);
when x"f3a" => lut_sig <= to_unsigned(integer(my_rom(3898)),16);
when x"f3b" => lut_sig <= to_unsigned(integer(my_rom(3899)),16);
when x"f3c" => lut_sig <= to_unsigned(integer(my_rom(3900)),16);
when x"f3d" => lut_sig <= to_unsigned(integer(my_rom(3901)),16);
when x"f3e" => lut_sig <= to_unsigned(integer(my_rom(3902)),16);
when x"f3f" => lut_sig <= to_unsigned(integer(my_rom(3903)),16);
when x"f40" => lut_sig <= to_unsigned(integer(my_rom(3904)),16);
when x"f41" => lut_sig <= to_unsigned(integer(my_rom(3905)),16);
when x"f42" => lut_sig <= to_unsigned(integer(my_rom(3906)),16);
when x"f43" => lut_sig <= to_unsigned(integer(my_rom(3907)),16);
when x"f44" => lut_sig <= to_unsigned(integer(my_rom(3908)),16);
when x"f45" => lut_sig <= to_unsigned(integer(my_rom(3909)),16);
when x"f46" => lut_sig <= to_unsigned(integer(my_rom(3910)),16);
when x"f47" => lut_sig <= to_unsigned(integer(my_rom(3911)),16);
when x"f48" => lut_sig <= to_unsigned(integer(my_rom(3912)),16);
when x"f49" => lut_sig <= to_unsigned(integer(my_rom(3913)),16);
when x"f4a" => lut_sig <= to_unsigned(integer(my_rom(3914)),16);
when x"f4b" => lut_sig <= to_unsigned(integer(my_rom(3915)),16);
when x"f4c" => lut_sig <= to_unsigned(integer(my_rom(3916)),16);
when x"f4d" => lut_sig <= to_unsigned(integer(my_rom(3917)),16);
when x"f4e" => lut_sig <= to_unsigned(integer(my_rom(3918)),16);
when x"f4f" => lut_sig <= to_unsigned(integer(my_rom(3919)),16);
when x"f50" => lut_sig <= to_unsigned(integer(my_rom(3920)),16);
when x"f51" => lut_sig <= to_unsigned(integer(my_rom(3921)),16);
when x"f52" => lut_sig <= to_unsigned(integer(my_rom(3922)),16);
when x"f53" => lut_sig <= to_unsigned(integer(my_rom(3923)),16);
when x"f54" => lut_sig <= to_unsigned(integer(my_rom(3924)),16);
when x"f55" => lut_sig <= to_unsigned(integer(my_rom(3925)),16);
when x"f56" => lut_sig <= to_unsigned(integer(my_rom(3926)),16);
when x"f57" => lut_sig <= to_unsigned(integer(my_rom(3927)),16);
when x"f58" => lut_sig <= to_unsigned(integer(my_rom(3928)),16);
when x"f59" => lut_sig <= to_unsigned(integer(my_rom(3929)),16);
when x"f5a" => lut_sig <= to_unsigned(integer(my_rom(3930)),16);
when x"f5b" => lut_sig <= to_unsigned(integer(my_rom(3931)),16);
when x"f5c" => lut_sig <= to_unsigned(integer(my_rom(3932)),16);
when x"f5d" => lut_sig <= to_unsigned(integer(my_rom(3933)),16);
when x"f5e" => lut_sig <= to_unsigned(integer(my_rom(3934)),16);
when x"f5f" => lut_sig <= to_unsigned(integer(my_rom(3935)),16);
when x"f60" => lut_sig <= to_unsigned(integer(my_rom(3936)),16);
when x"f61" => lut_sig <= to_unsigned(integer(my_rom(3937)),16);
when x"f62" => lut_sig <= to_unsigned(integer(my_rom(3938)),16);
when x"f63" => lut_sig <= to_unsigned(integer(my_rom(3939)),16);
when x"f64" => lut_sig <= to_unsigned(integer(my_rom(3940)),16);
when x"f65" => lut_sig <= to_unsigned(integer(my_rom(3941)),16);
when x"f66" => lut_sig <= to_unsigned(integer(my_rom(3942)),16);
when x"f67" => lut_sig <= to_unsigned(integer(my_rom(3943)),16);
when x"f68" => lut_sig <= to_unsigned(integer(my_rom(3944)),16);
when x"f69" => lut_sig <= to_unsigned(integer(my_rom(3945)),16);
when x"f6a" => lut_sig <= to_unsigned(integer(my_rom(3946)),16);
when x"f6b" => lut_sig <= to_unsigned(integer(my_rom(3947)),16);
when x"f6c" => lut_sig <= to_unsigned(integer(my_rom(3948)),16);
when x"f6d" => lut_sig <= to_unsigned(integer(my_rom(3949)),16);
when x"f6e" => lut_sig <= to_unsigned(integer(my_rom(3950)),16);
when x"f6f" => lut_sig <= to_unsigned(integer(my_rom(3951)),16);
when x"f70" => lut_sig <= to_unsigned(integer(my_rom(3952)),16);
when x"f71" => lut_sig <= to_unsigned(integer(my_rom(3953)),16);
when x"f72" => lut_sig <= to_unsigned(integer(my_rom(3954)),16);
when x"f73" => lut_sig <= to_unsigned(integer(my_rom(3955)),16);
when x"f74" => lut_sig <= to_unsigned(integer(my_rom(3956)),16);
when x"f75" => lut_sig <= to_unsigned(integer(my_rom(3957)),16);
when x"f76" => lut_sig <= to_unsigned(integer(my_rom(3958)),16);
when x"f77" => lut_sig <= to_unsigned(integer(my_rom(3959)),16);
when x"f78" => lut_sig <= to_unsigned(integer(my_rom(3960)),16);
when x"f79" => lut_sig <= to_unsigned(integer(my_rom(3961)),16);
when x"f7a" => lut_sig <= to_unsigned(integer(my_rom(3962)),16);
when x"f7b" => lut_sig <= to_unsigned(integer(my_rom(3963)),16);
when x"f7c" => lut_sig <= to_unsigned(integer(my_rom(3964)),16);
when x"f7d" => lut_sig <= to_unsigned(integer(my_rom(3965)),16);
when x"f7e" => lut_sig <= to_unsigned(integer(my_rom(3966)),16);
when x"f7f" => lut_sig <= to_unsigned(integer(my_rom(3967)),16);
when x"f80" => lut_sig <= to_unsigned(integer(my_rom(3968)),16);
when x"f81" => lut_sig <= to_unsigned(integer(my_rom(3969)),16);
when x"f82" => lut_sig <= to_unsigned(integer(my_rom(3970)),16);
when x"f83" => lut_sig <= to_unsigned(integer(my_rom(3971)),16);
when x"f84" => lut_sig <= to_unsigned(integer(my_rom(3972)),16);
when x"f85" => lut_sig <= to_unsigned(integer(my_rom(3973)),16);
when x"f86" => lut_sig <= to_unsigned(integer(my_rom(3974)),16);
when x"f87" => lut_sig <= to_unsigned(integer(my_rom(3975)),16);
when x"f88" => lut_sig <= to_unsigned(integer(my_rom(3976)),16);
when x"f89" => lut_sig <= to_unsigned(integer(my_rom(3977)),16);
when x"f8a" => lut_sig <= to_unsigned(integer(my_rom(3978)),16);
when x"f8b" => lut_sig <= to_unsigned(integer(my_rom(3979)),16);
when x"f8c" => lut_sig <= to_unsigned(integer(my_rom(3980)),16);
when x"f8d" => lut_sig <= to_unsigned(integer(my_rom(3981)),16);
when x"f8e" => lut_sig <= to_unsigned(integer(my_rom(3982)),16);
when x"f8f" => lut_sig <= to_unsigned(integer(my_rom(3983)),16);
when x"f90" => lut_sig <= to_unsigned(integer(my_rom(3984)),16);
when x"f91" => lut_sig <= to_unsigned(integer(my_rom(3985)),16);
when x"f92" => lut_sig <= to_unsigned(integer(my_rom(3986)),16);
when x"f93" => lut_sig <= to_unsigned(integer(my_rom(3987)),16);
when x"f94" => lut_sig <= to_unsigned(integer(my_rom(3988)),16);
when x"f95" => lut_sig <= to_unsigned(integer(my_rom(3989)),16);
when x"f96" => lut_sig <= to_unsigned(integer(my_rom(3990)),16);
when x"f97" => lut_sig <= to_unsigned(integer(my_rom(3991)),16);
when x"f98" => lut_sig <= to_unsigned(integer(my_rom(3992)),16);
when x"f99" => lut_sig <= to_unsigned(integer(my_rom(3993)),16);
when x"f9a" => lut_sig <= to_unsigned(integer(my_rom(3994)),16);
when x"f9b" => lut_sig <= to_unsigned(integer(my_rom(3995)),16);
when x"f9c" => lut_sig <= to_unsigned(integer(my_rom(3996)),16);
when x"f9d" => lut_sig <= to_unsigned(integer(my_rom(3997)),16);
when x"f9e" => lut_sig <= to_unsigned(integer(my_rom(3998)),16);
when x"f9f" => lut_sig <= to_unsigned(integer(my_rom(3999)),16);
when x"fa0" => lut_sig <= to_unsigned(integer(my_rom(4000)),16);
when x"fa1" => lut_sig <= to_unsigned(integer(my_rom(4001)),16);
when x"fa2" => lut_sig <= to_unsigned(integer(my_rom(4002)),16);
when x"fa3" => lut_sig <= to_unsigned(integer(my_rom(4003)),16);
when x"fa4" => lut_sig <= to_unsigned(integer(my_rom(4004)),16);
when x"fa5" => lut_sig <= to_unsigned(integer(my_rom(4005)),16);
when x"fa6" => lut_sig <= to_unsigned(integer(my_rom(4006)),16);
when x"fa7" => lut_sig <= to_unsigned(integer(my_rom(4007)),16);
when x"fa8" => lut_sig <= to_unsigned(integer(my_rom(4008)),16);
when x"fa9" => lut_sig <= to_unsigned(integer(my_rom(4009)),16);
when x"faa" => lut_sig <= to_unsigned(integer(my_rom(4010)),16);
when x"fab" => lut_sig <= to_unsigned(integer(my_rom(4011)),16);
when x"fac" => lut_sig <= to_unsigned(integer(my_rom(4012)),16);
when x"fad" => lut_sig <= to_unsigned(integer(my_rom(4013)),16);
when x"fae" => lut_sig <= to_unsigned(integer(my_rom(4014)),16);
when x"faf" => lut_sig <= to_unsigned(integer(my_rom(4015)),16);
when x"fb0" => lut_sig <= to_unsigned(integer(my_rom(4016)),16);
when x"fb1" => lut_sig <= to_unsigned(integer(my_rom(4017)),16);
when x"fb2" => lut_sig <= to_unsigned(integer(my_rom(4018)),16);
when x"fb3" => lut_sig <= to_unsigned(integer(my_rom(4019)),16);
when x"fb4" => lut_sig <= to_unsigned(integer(my_rom(4020)),16);
when x"fb5" => lut_sig <= to_unsigned(integer(my_rom(4021)),16);
when x"fb6" => lut_sig <= to_unsigned(integer(my_rom(4022)),16);
when x"fb7" => lut_sig <= to_unsigned(integer(my_rom(4023)),16);
when x"fb8" => lut_sig <= to_unsigned(integer(my_rom(4024)),16);
when x"fb9" => lut_sig <= to_unsigned(integer(my_rom(4025)),16);
when x"fba" => lut_sig <= to_unsigned(integer(my_rom(4026)),16);
when x"fbb" => lut_sig <= to_unsigned(integer(my_rom(4027)),16);
when x"fbc" => lut_sig <= to_unsigned(integer(my_rom(4028)),16);
when x"fbd" => lut_sig <= to_unsigned(integer(my_rom(4029)),16);
when x"fbe" => lut_sig <= to_unsigned(integer(my_rom(4030)),16);
when x"fbf" => lut_sig <= to_unsigned(integer(my_rom(4031)),16);
when x"fc0" => lut_sig <= to_unsigned(integer(my_rom(4032)),16);
when x"fc1" => lut_sig <= to_unsigned(integer(my_rom(4033)),16);
when x"fc2" => lut_sig <= to_unsigned(integer(my_rom(4034)),16);
when x"fc3" => lut_sig <= to_unsigned(integer(my_rom(4035)),16);
when x"fc4" => lut_sig <= to_unsigned(integer(my_rom(4036)),16);
when x"fc5" => lut_sig <= to_unsigned(integer(my_rom(4037)),16);
when x"fc6" => lut_sig <= to_unsigned(integer(my_rom(4038)),16);
when x"fc7" => lut_sig <= to_unsigned(integer(my_rom(4039)),16);
when x"fc8" => lut_sig <= to_unsigned(integer(my_rom(4040)),16);
when x"fc9" => lut_sig <= to_unsigned(integer(my_rom(4041)),16);
when x"fca" => lut_sig <= to_unsigned(integer(my_rom(4042)),16);
when x"fcb" => lut_sig <= to_unsigned(integer(my_rom(4043)),16);
when x"fcc" => lut_sig <= to_unsigned(integer(my_rom(4044)),16);
when x"fcd" => lut_sig <= to_unsigned(integer(my_rom(4045)),16);
when x"fce" => lut_sig <= to_unsigned(integer(my_rom(4046)),16);
when x"fcf" => lut_sig <= to_unsigned(integer(my_rom(4047)),16);
when x"fd0" => lut_sig <= to_unsigned(integer(my_rom(4048)),16);
when x"fd1" => lut_sig <= to_unsigned(integer(my_rom(4049)),16);
when x"fd2" => lut_sig <= to_unsigned(integer(my_rom(4050)),16);
when x"fd3" => lut_sig <= to_unsigned(integer(my_rom(4051)),16);
when x"fd4" => lut_sig <= to_unsigned(integer(my_rom(4052)),16);
when x"fd5" => lut_sig <= to_unsigned(integer(my_rom(4053)),16);
when x"fd6" => lut_sig <= to_unsigned(integer(my_rom(4054)),16);
when x"fd7" => lut_sig <= to_unsigned(integer(my_rom(4055)),16);
when x"fd8" => lut_sig <= to_unsigned(integer(my_rom(4056)),16);
when x"fd9" => lut_sig <= to_unsigned(integer(my_rom(4057)),16);
when x"fda" => lut_sig <= to_unsigned(integer(my_rom(4058)),16);
when x"fdb" => lut_sig <= to_unsigned(integer(my_rom(4059)),16);
when x"fdc" => lut_sig <= to_unsigned(integer(my_rom(4060)),16);
when x"fdd" => lut_sig <= to_unsigned(integer(my_rom(4061)),16);
when x"fde" => lut_sig <= to_unsigned(integer(my_rom(4062)),16);
when x"fdf" => lut_sig <= to_unsigned(integer(my_rom(4063)),16);
when x"fe0" => lut_sig <= to_unsigned(integer(my_rom(4064)),16);
when x"fe1" => lut_sig <= to_unsigned(integer(my_rom(4065)),16);
when x"fe2" => lut_sig <= to_unsigned(integer(my_rom(4066)),16);
when x"fe3" => lut_sig <= to_unsigned(integer(my_rom(4067)),16);
when x"fe4" => lut_sig <= to_unsigned(integer(my_rom(4068)),16);
when x"fe5" => lut_sig <= to_unsigned(integer(my_rom(4069)),16);
when x"fe6" => lut_sig <= to_unsigned(integer(my_rom(4070)),16);
when x"fe7" => lut_sig <= to_unsigned(integer(my_rom(4071)),16);
when x"fe8" => lut_sig <= to_unsigned(integer(my_rom(4072)),16);
when x"fe9" => lut_sig <= to_unsigned(integer(my_rom(4073)),16);
when x"fea" => lut_sig <= to_unsigned(integer(my_rom(4074)),16);
when x"feb" => lut_sig <= to_unsigned(integer(my_rom(4075)),16);
when x"fec" => lut_sig <= to_unsigned(integer(my_rom(4076)),16);
when x"fed" => lut_sig <= to_unsigned(integer(my_rom(4077)),16);
when x"fee" => lut_sig <= to_unsigned(integer(my_rom(4078)),16);
when x"fef" => lut_sig <= to_unsigned(integer(my_rom(4079)),16);
when x"ff0" => lut_sig <= to_unsigned(integer(my_rom(4080)),16);
when x"ff1" => lut_sig <= to_unsigned(integer(my_rom(4081)),16);
when x"ff2" => lut_sig <= to_unsigned(integer(my_rom(4082)),16);
when x"ff3" => lut_sig <= to_unsigned(integer(my_rom(4083)),16);
when x"ff4" => lut_sig <= to_unsigned(integer(my_rom(4084)),16);
when x"ff5" => lut_sig <= to_unsigned(integer(my_rom(4085)),16);
when x"ff6" => lut_sig <= to_unsigned(integer(my_rom(4086)),16);
when x"ff7" => lut_sig <= to_unsigned(integer(my_rom(4087)),16);
when x"ff8" => lut_sig <= to_unsigned(integer(my_rom(4088)),16);
when x"ff9" => lut_sig <= to_unsigned(integer(my_rom(4089)),16);
when x"ffa" => lut_sig <= to_unsigned(integer(my_rom(4090)),16);
when x"ffb" => lut_sig <= to_unsigned(integer(my_rom(4091)),16);
when x"ffc" => lut_sig <= to_unsigned(integer(my_rom(4092)),16);
when x"ffd" => lut_sig <= to_unsigned(integer(my_rom(4093)),16);
when x"ffe" => lut_sig <= to_unsigned(integer(my_rom(4094)),16);
when x"fff" => lut_sig <= to_unsigned(integer(my_rom(4095)),16);
                    when others => lut_sig <= "0000000000000000";
                end case;
            end process;
end Behavioral;
