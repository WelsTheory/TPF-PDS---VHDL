library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cos_entity is
    Port (
        address: in std_logic_vector(11 downto 0);
        cos: out std_logic_vector(15 downto 0)
    );
end entity;

architecture Behavioral of cos_entity is
    
    type mem is array(0 to 4095) of real;
    constant my_cos: mem := (
0=>1500.0,
1=>1499.999117157754,
2=>1499.9964686330936,
3=>1499.992054432255,
4=>1499.9858745656297,
5=>1499.9779290477668,
6=>1499.9682178973721,
7=>1499.9567411373077,
8=>1499.9434987945933,
9=>1499.928490900404,
10=>1499.9117174900723,
11=>1499.893178603087,
12=>1499.8728742830936,
13=>1499.8508045778926,
14=>1499.8269695394422,
15=>1499.8013692238555,
16=>1499.7740036914024,
17=>1499.7448730065078,
18=>1499.7139772377525,
19=>1499.6813164578728,
20=>1499.6468907437602,
21=>1499.6107001764613,
22=>1499.5727448411776,
23=>1499.5330248272653,
24=>1499.491540228235,
25=>1499.4482911417517,
26=>1499.4032776696345,
27=>1499.3564999178561,
28=>1499.3079579965429,
29=>1499.257652019974,
30=>1499.205582106583,
31=>1499.1517483789548,
32=>1499.0961509638269,
33=>1499.0387899920897,
34=>1498.9796655987852,
35=>1498.9187779231063,
36=>1498.856127108398,
37=>1498.7917133021551,
38=>1498.7255366560244,
39=>1498.6575973258014,
40=>1498.5878954714321,
41=>1498.5164312570118,
42=>1498.4432048507852,
43=>1498.3682164251447,
44=>1498.291466156632,
45=>1498.2129542259358,
46=>1498.1326808178924,
47=>1498.0506461214854,
48=>1497.9668503298449,
49=>1497.8812936402464,
50=>1497.7939762541114,
51=>1497.7048983770064,
52=>1497.6140602186433,
53=>1497.5214619928765,
54=>1497.427103917706,
55=>1497.3309862152732,
56=>1497.233109111863,
57=>1497.1334728379022,
58=>1497.032077627959,
59=>1496.9289237207431,
60=>1496.824011359104,
61=>1496.7173407900307,
62=>1496.6089122646524,
63=>1496.4987260382363,
64=>1496.3867823701885,
65=>1496.2730815240511,
66=>1496.1576237675042,
67=>1496.040409372364,
68=>1495.9214386145816,
69=>1495.8007117742436,
70=>1495.6782291355707,
71=>1495.5539909869176,
72=>1495.4279976207708,
73=>1495.30024933375,
74=>1495.1707464266055,
75=>1495.03948920422,
76=>1494.9064779756045,
77=>1494.7717130539008,
78=>1494.635194756378,
79=>1494.4969234044343,
80=>1494.356899323594,
81=>1494.2151228435087,
82=>1494.0715942979548,
83=>1493.926314024834,
84=>1493.7792823661716,
85=>1493.6304996681163,
86=>1493.4799662809394,
87=>1493.3276825590333,
88=>1493.1736488609115,
89=>1493.0178655492073,
90=>1492.8603329906723,
91=>1492.7010515561778,
92=>1492.5400216207108,
93=>1492.3772435633757,
94=>1492.2127177673922,
95=>1492.046444620094,
96=>1491.8784245129295,
97=>1491.7086578414592,
98=>1491.5371450053553,
99=>1491.3638864084019,
100=>1491.1888824584917,
101=>1491.0121335676274,
102=>1490.833640151919,
103=>1490.6534026315844,
104=>1490.4714214309467,
105=>1490.2876969784347,
106=>1490.1022297065806,
107=>1489.9150200520203,
108=>1489.7260684554913,
109=>1489.5353753618317,
110=>1489.3429412199807,
111=>1489.1487664829751,
112=>1488.9528516079502,
113=>1488.7551970561376,
114=>1488.555803292865,
115=>1488.3546707875544,
116=>1488.1518000137207,
117=>1487.9471914489723,
118=>1487.7408455750076,
119=>1487.5327628776156,
120=>1487.3229438466742,
121=>1487.1113889761493,
122=>1486.8980987640928,
123=>1486.6830737126422,
124=>1486.4663143280197,
125=>1486.24782112053,
126=>1486.02759460456,
127=>1485.805635298577,
128=>1485.581943725128,
129=>1485.3565204108377,
130=>1485.1293658864079,
131=>1484.9004806866164,
132=>1484.6698653503158,
133=>1484.4375204204307,
134=>1484.2034464439585,
135=>1483.9676439719665,
136=>1483.7301135595922,
137=>1483.4908557660403,
138=>1483.2498711545827,
139=>1483.0071602925568,
140=>1482.762723751363,
141=>1482.5165621064652,
142=>1482.2686759373887,
143=>1482.0190658277184,
144=>1481.7677323650978,
145=>1481.514676141228,
146=>1481.2598977518653,
147=>1481.003397796821,
148=>1480.7451768799588,
149=>1480.4852356091942,
150=>1480.223574596493,
151=>1479.9601944578699,
152=>1479.6950958133862,
153=>1479.4282792871495,
154=>1479.1597455073115,
155=>1478.8894951060665,
156=>1478.6175287196506,
157=>1478.3438469883397,
158=>1478.0684505564477,
159=>1477.791340072326,
160=>1477.5125161883602,
161=>1477.2319795609708,
162=>1476.9497308506097,
163=>1476.66577072176,
164=>1476.3800998429338,
165=>1476.0927188866704,
166=>1475.8036285295352,
167=>1475.5128294521185,
168=>1475.2203223390322,
169=>1474.9261078789104,
170=>1474.630186764406,
171=>1474.332559692191,
172=>1474.0332273629513,
173=>1473.7321904813898,
174=>1473.4294497562214,
175=>1473.1250059001718,
176=>1472.818859629977,
177=>1472.5110116663805,
178=>1472.2014627341323,
179=>1471.8902135619865,
180=>1471.5772648827005,
181=>1471.2626174330321,
182=>1470.9462719537391,
183=>1470.6282291895766,
184=>1470.3084898892953,
185=>1469.9870548056401,
186=>1469.6639246953487,
187=>1469.3391003191487,
188=>1469.012582441756,
189=>1468.6843718318746,
190=>1468.354469262193,
191=>1468.0228755093829,
192=>1467.6895913540975,
193=>1467.3546175809697,
194=>1467.0179549786103,
195=>1466.6796043396057,
196=>1466.3395664605164,
197=>1465.9978421418755,
198=>1465.654432188186,
199=>1465.3093374079199,
200=>1464.9625586135144,
201=>1464.6140966213725,
202=>1464.2639522518593,
203=>1463.912126329301,
204=>1463.5586196819818,
205=>1463.2034331421441,
206=>1462.8465675459838,
207=>1462.4880237336506,
208=>1462.1278025492447,
209=>1461.7659048408154,
210=>1461.4023314603592,
211=>1461.0370832638168,
212=>1460.6701611110725,
213=>1460.3015658659515,
214=>1459.9312983962172,
215=>1459.5593595735709,
216=>1459.1857502736477,
217=>1458.810471376016,
218=>1458.4335237641744,
219=>1458.0549083255505,
220=>1457.674625951498,
221=>1457.2926775372953,
222=>1456.909063982143,
223=>1456.5237861891615,
224=>1456.13684506539,
225=>1455.7482415217823,
226=>1455.3579764732076,
227=>1454.966050838445,
228=>1454.5724655401846,
229=>1454.1772215050223,
230=>1453.7803196634604,
231=>1453.3817609499033,
232=>1452.9815463026562,
233=>1452.5796766639228,
234=>1452.1761529798027,
235=>1451.7709762002908,
236=>1451.3641472792724,
237=>1450.9556671745227,
238=>1450.5455368477046,
239=>1450.1337572643656,
240=>1449.720329393936,
241=>1449.3052542097275,
242=>1448.8885326889283,
243=>1448.4701658126037,
244=>1448.050154565692,
245=>1447.6284999370037,
246=>1447.2052029192168,
247=>1446.7802645088768,
248=>1446.3536857063937,
249=>1445.9254675160382,
250=>1445.4956109459417,
251=>1445.0641170080921,
252=>1444.6309867183322,
253=>1444.196221096358,
254=>1443.7598211657137,
255=>1443.3217879537924,
256=>1442.8821224918324,
257=>1442.4408258149142,
258=>1441.9978989619585,
259=>1441.5533429757243,
260=>1441.1071589028056,
261=>1440.6593477936296,
262=>1440.2099107024537,
263=>1439.7588486873635,
264=>1439.3061628102698,
265=>1438.8518541369065,
266=>1438.395923736828,
267=>1437.9383726834067,
268=>1437.4792020538302,
269=>1437.0184129290992,
270=>1436.5560063940247,
271=>1436.0919835372254,
272=>1435.6263454511252,
273=>1435.1590932319507,
274=>1434.6902279797287,
275=>1434.2197507982828,
276=>1433.7476627952328,
277=>1433.2739650819897,
278=>1432.7986587737541,
279=>1432.3217449895144,
280=>1431.8432248520428,
281=>1431.3630994878934,
282=>1430.8813700273995,
283=>1430.3980376046704,
284=>1429.91310335759,
285=>1429.4265684278125,
286=>1428.938433960761,
287=>1428.448701105624,
288=>1427.9573710153531,
289=>1427.4644448466606,
290=>1426.9699237600153,
291=>1426.4738089196417,
292=>1425.9761014935161,
293=>1425.4768026533645,
294=>1424.975913574659,
295=>1424.473435436616,
296=>1423.9693694221924,
297=>1423.463716718083,
298=>1422.9564785147197,
299=>1422.4476560062656,
300=>1421.9372503906138,
301=>1421.425262869385,
302=>1420.9116946479235,
303=>1420.3965469352956,
304=>1419.8798209442853,
305=>1419.3615178913929,
306=>1418.8416389968315,
307=>1418.3201854845233,
308=>1417.7971585820987,
309=>1417.2725595208917,
310=>1416.746389535937,
311=>1416.2186498659687,
312=>1415.6893417534156,
313=>1415.1584664443992,
314=>1414.6260251887306,
315=>1414.0920192399076,
316=>1413.5564498551112,
317=>1413.019318295204,
318=>1412.4806258247252,
319=>1411.9403737118898,
320=>1411.3985632285844,
321=>1410.8551956503634,
322=>1410.3102722564486,
323=>1409.7637943297232,
324=>1409.2157631567306,
325=>1408.6661800276715,
326=>1408.1150462363992,
327=>1407.5623630804184,
328=>1407.0081318608816,
329=>1406.4523538825847,
330=>1405.8950304539667,
331=>1405.336162887103,
332=>1404.775752497706,
333=>1404.2138006051196,
334=>1403.6503085323166,
335=>1403.085277605896,
336=>1402.5187091560795,
337=>1401.9506045167086,
338=>1401.3809650252417,
339=>1400.8097920227501,
340=>1400.2370868539151,
341=>1399.6628508670265,
342=>1399.0870854139762,
343=>1398.509791850258,
344=>1397.9309715349632,
345=>1397.3506258307766,
346=>1396.7687561039756,
347=>1396.185363724424,
348=>1395.600450065571,
349=>1395.0140165044477,
350=>1394.4260644216627,
351=>1393.8365952013996,
352=>1393.2456102314143,
353=>1392.6531109030307,
354=>1392.0590986111376,
355=>1391.4635747541865,
356=>1390.8665407341873,
357=>1390.2679979567042,
358=>1389.6679478308547,
359=>1389.0663917693041,
360=>1388.4633311882635,
361=>1387.8587675074857,
362=>1387.2527021502624,
363=>1386.645136543421,
364=>1386.0360721173195,
365=>1385.425510305846,
366=>1384.813452546413,
367=>1384.1999002799553,
368=>1383.5848549509253,
369=>1382.9683180072916,
370=>1382.3502909005333,
371=>1381.7307750856387,
372=>1381.1097720211,
373=>1380.4872831689117,
374=>1379.863309994565,
375=>1379.237853967047,
376=>1378.6109165588346,
377=>1377.9824992458925,
378=>1377.3526035076702,
379=>1376.7212308270964,
380=>1376.0883826905788,
381=>1375.4540605879965,
382=>1374.8182660127006,
383=>1374.1810004615074,
384=>1373.5422654346971,
385=>1372.9020624360087,
386=>1372.2603929726379,
387=>1371.6172585552324,
388=>1370.9726606978886,
389=>1370.3266009181486,
390=>1369.6790807369962,
391=>1369.0301016788528,
392=>1368.379665271575,
393=>1367.7277730464502,
394=>1367.0744265381927,
395=>1366.4196272849413,
396=>1365.763376828254,
397=>1365.1056767131065,
398=>1364.446528487886,
399=>1363.7859337043901,
400=>1363.123893917821,
401=>1362.4604106867837,
402=>1361.7954855732805,
403=>1361.1291201427089,
404=>1360.4613159638566,
405=>1359.7920746088994,
406=>1359.121397653396,
407=>1358.4492866762848,
408=>1357.7757432598805,
409=>1357.1007689898697,
410=>1356.4243654553084,
411=>1355.7465342486166,
412=>1355.0672769655757,
413=>1354.3865952053243,
414=>1353.704490570355,
415=>1353.0209646665094,
416=>1352.3360191029765,
417=>1351.6496554922855,
418=>1350.9618754503063,
419=>1350.2726805962416,
420=>1349.582072552626,
421=>1348.8900529453203,
422=>1348.1966234035092,
423=>1347.5017855596961,
424=>1346.8055410497009,
425=>1346.1078915126536,
426=>1345.4088385909936,
427=>1344.7083839304628,
428=>1344.0065291801038,
429=>1343.303275992256,
430=>1342.5986260225498,
431=>1341.8925809299046,
432=>1341.1851423765243,
433=>1340.4763120278935,
434=>1339.766091552773,
435=>1339.0544826231967,
436=>1338.3414869144667,
437=>1337.6271061051507,
438=>1336.9113418770762,
439=>1336.1941959153291,
440=>1335.4756699082468,
441=>1334.7557655474168,
442=>1334.0344845276704,
443=>1333.3118285470812,
444=>1332.587799306959,
445=>1331.862398511846,
446=>1331.1356278695148,
447=>1330.4074890909624,
448=>1329.6779838904063,
449=>1328.9471139852812,
450=>1328.2148810962346,
451=>1327.4812869471232,
452=>1326.7463332650077,
453=>1326.0100217801498,
454=>1325.2723542260082,
455=>1324.5333323392335,
456=>1323.7929578596654,
457=>1323.051232530327,
458=>1322.3081580974224,
459=>1321.563736310332,
460=>1320.8179689216072,
461=>1320.0708576869683,
462=>1319.3224043652986,
463=>1318.5726107186417,
464=>1317.821478512196,
465=>1317.0690095143118,
466=>1316.3152054964858,
467=>1315.5600682333584,
468=>1314.8035995027083,
469=>1314.045801085449,
470=>1313.2866747656244,
471=>1312.5262223304048,
472=>1311.764445570082,
473=>1311.001346278066,
474=>1310.2369262508803,
475=>1309.4711872881576,
476=>1308.7041311926357,
477=>1307.9357597701537,
478=>1307.1660748296465,
479=>1306.395078183142,
480=>1305.622771645756,
481=>1304.849157035688,
482=>1304.0742361742173,
483=>1303.2980108856977,
484=>1302.5204829975548,
485=>1301.7416543402808,
486=>1300.9615267474294,
487=>1300.1801020556131,
488=>1299.3973821044983,
489=>1298.6133687367992,
490=>1297.8280637982775,
491=>1297.041469137733,
492=>1296.2535866070036,
493=>1295.4644180609587,
494=>1294.673965357495,
495=>1293.8822303575325,
496=>1293.08921492501,
497=>1292.2949209268816,
498=>1291.4993502331101,
499=>1290.7025047166649,
500=>1289.9043862535163,
501=>1289.1049967226313,
502=>1288.3043380059698,
503=>1287.5024119884793,
504=>1286.6992205580907,
505=>1285.8947656057146,
506=>1285.0890490252355,
507=>1284.2820727135086,
508=>1283.4738385703545,
509=>1282.6643484985552,
510=>1281.8536044038499,
511=>1281.0416081949288,
512=>1280.2283617834316,
513=>1279.4138670839397,
514=>1278.5981260139747,
515=>1277.7811404939907,
516=>1276.9629124473736,
517=>1276.143443800433,
518=>1275.3227364823997,
519=>1274.500792425421,
520=>1273.6776135645546,
521=>1272.8532018377668,
522=>1272.0275591859254,
523=>1271.200687552796,
524=>1270.372588885038,
525=>1269.5432651321996,
526=>1268.7127182467125,
527=>1267.880950183889,
528=>1267.047962901915,
529=>1266.2137583618478,
530=>1265.3783385276101,
531=>1264.541705365986,
532=>1263.703860846615,
533=>1262.86480694199,
534=>1262.02454562745,
535=>1261.1830788811765,
536=>1260.3404086841897,
537=>1259.4965370203422,
538=>1258.6514658763156,
539=>1257.8051972416154,
540=>1256.9577331085657,
541=>1256.1090754723061,
542=>1255.259226330785,
543=>1254.4081876847565,
544=>1253.5559615377751,
545=>1252.7025498961905,
546=>1251.8479547691436,
547=>1250.9921781685618,
548=>1250.1352221091538,
549=>1249.2770886084045,
550=>1248.4177796865717,
551=>1247.55729736668,
552=>1246.6956436745158,
553=>1245.8328206386248,
554=>1244.968830290304,
555=>1244.1036746635993,
556=>1243.2373557953001,
557=>1242.369875724934,
558=>1241.5012364947625,
559=>1240.631440149776,
560=>1239.7604887376888,
561=>1238.8883843089352,
562=>1238.0151289166636,
563=>1237.1407246167314,
564=>1236.265173467702,
565=>1235.388477530838,
566=>1234.5106388700972,
567=>1233.631659552128,
568=>1232.7515416462636,
569=>1231.870287224518,
570=>1230.9878983615818,
571=>1230.104377134814,
572=>1229.219725624242,
573=>1228.3339459125525,
574=>1227.4470400850892,
575=>1226.5590102298463,
576=>1225.6698584374649,
577=>1224.7795868012267,
578=>1223.8881974170502,
579=>1222.9956923834852,
580=>1222.1020738017085,
581=>1221.2073437755175,
582=>1220.3115044113272,
583=>1219.4145578181635,
584=>1218.5165061076598,
585=>1217.6173513940503,
586=>1216.7170957941664,
587=>1215.8157414274315,
588=>1214.9132904158553,
589=>1214.0097448840295,
590=>1213.1051069591226,
591=>1212.1993787708748,
592=>1211.292562451593,
593=>1210.3846601361458,
594=>1209.4756739619588,
595=>1208.5656060690092,
596=>1207.6544585998201,
597=>1206.7422336994573,
598=>1205.8289335155225,
599=>1204.9145601981488,
600=>1203.999115899996,
601=>1203.0826027762455,
602=>1202.165022984594,
603=>1201.2463786852509,
604=>1200.32667204093,
605=>1199.4059052168473,
606=>1198.4840803807144,
607=>1197.561199702734,
608=>1196.637265355594,
609=>1195.7122795144633,
610=>1194.7862443569857,
611=>1193.8591620632758,
612=>1192.9310348159138,
613=>1192.0018647999395,
614=>1191.0716542028472,
615=>1190.140405214582,
616=>1189.2081200275327,
617=>1188.2748008365284,
618=>1187.3404498388313,
619=>1186.4050692341343,
620=>1185.4686612245532,
621=>1184.5312280146227,
622=>1183.5927718112912,
623=>1182.6532948239153,
624=>1181.7127992642552,
625=>1180.7712873464686,
626=>1179.8287612871063,
627=>1178.8852233051064,
628=>1177.9406756217895,
629=>1176.9951204608533,
630=>1176.0485600483669,
631=>1175.1009966127665,
632=>1174.1524323848496,
633=>1173.2028695977697,
634=>1172.2523104870313,
635=>1171.3007572904842,
636=>1170.3482122483188,
637=>1169.39467760306,
638=>1168.4401555995637,
639=>1167.484648485009,
640=>1166.5281585088949,
641=>1165.5706879230338,
642=>1164.6122389815473,
643=>1163.6528139408597,
644=>1162.692415059694,
645=>1161.731044599065,
646=>1160.7687048222754,
647=>1159.8053979949095,
648=>1158.8411263848288,
649=>1157.8758922621662,
650=>1156.9096978993196,
651=>1155.9425455709486,
652=>1154.9744375539676,
653=>1154.005376127541,
654=>1153.0353635730776,
655=>1152.0644021742262,
656=>1151.092494216868,
657=>1150.1196419891137,
658=>1149.145847781297,
659=>1148.1711138859687,
660=>1147.1954425978925,
661=>1146.2188362140382,
662=>1145.2412970335777,
663=>1144.2628273578785,
664=>1143.2834294904992,
665=>1142.3031057371832,
666=>1141.3218584058536,
667=>1140.3396898066082,
668=>1139.3566022517136,
669=>1138.3725980555994,
670=>1137.3876795348535,
671=>1136.401849008217,
672=>1135.4151087965765,
673=>1134.427461222962,
674=>1133.4389086125384,
675=>1132.449453292602,
676=>1131.4590975925737,
677=>1130.4678438439948,
678=>1129.4756943805203,
679=>1128.482651537914,
680=>1127.488717654043,
681=>1126.4938950688725,
682=>1125.4981861244592,
683=>1124.501593164947,
684=>1123.5041185365608,
685=>1122.5057645876018,
686=>1121.50653366844,
687=>1120.5064281315113,
688=>1119.5054503313097,
689=>1118.5036026243833,
690=>1117.5008873693287,
691=>1116.4973069267835,
692=>1115.4928636594234,
693=>1114.4875599319546,
694=>1113.4813981111095,
695=>1112.4743805656403,
696=>1111.4665096663146,
697=>1110.4577877859078,
698=>1109.4482172991998,
699=>1108.4378005829676,
700=>1107.426540015981,
701=>1106.4144379789957,
702=>1105.401496854749,
703=>1104.3877190279536,
704=>1103.3731068852921,
705=>1102.3576628154105,
706=>1101.3413892089143,
707=>1100.3242884583615,
708=>1099.3063629582575,
709=>1098.2876151050496,
710=>1097.2680472971201,
711=>1096.247661934783,
712=>1095.2264614202763,
713=>1094.2044481577573,
714=>1093.1816245532966,
715=>1092.1579930148723,
716=>1091.1335559523652,
717=>1090.108315777552,
718=>1089.0822749041004,
719=>1088.0554357475626,
720=>1087.027800725371,
721=>1085.999372256831,
722=>1084.9701527631164,
723=>1083.940144667263,
724=>1082.909350394163,
725=>1081.8777723705603,
726=>1080.8454130250425,
727=>1079.812274788038,
728=>1078.778360091808,
729=>1077.7436713704424,
730=>1076.7082110598528,
731=>1075.6719815977674,
732=>1074.6349854237253,
733=>1073.5972249790707,
734=>1072.5587027069469,
735=>1071.5194210522907,
736=>1070.4793824618268,
737=>1069.4385893840622,
738=>1068.3970442692791,
739=>1067.3547495695316,
740=>1066.3117077386376,
741=>1065.267921232174,
742=>1064.2233925074715,
743=>1063.1781240236069,
744=>1062.1321182414,
745=>1061.0853776234053,
746=>1060.0379046339076,
747=>1058.9897017389167,
748=>1057.9407714061592,
749=>1056.8911161050755,
750=>1055.8407383068127,
751=>1054.7896404842181,
752=>1053.7378251118346,
753=>1052.6852946658944,
754=>1051.6320516243131,
755=>1050.5780984666837,
756=>1049.5234376742715,
757=>1048.4680717300075,
758=>1047.4120031184823,
759=>1046.3552343259414,
760=>1045.2977678402788,
761=>1044.2396061510303,
762=>1043.180751749369,
763=>1042.1212071280986,
764=>1041.0609747816477,
765=>1040.0000572060642,
766=>1038.9384568990088,
767=>1037.8761763597504,
768=>1036.8132180891578,
769=>1035.7495845896967,
770=>1034.6852783654224,
771=>1033.620301921973,
772=>1032.5546577665648,
773=>1031.488348407987,
774=>1030.4213763565938,
775=>1029.3537441242997,
776=>1028.2854542245736,
777=>1027.2165091724332,
778=>1026.1469114844376,
779=>1025.0766636786832,
780=>1024.0057682747965,
781=>1022.9342277939284,
782=>1021.8620447587491,
783=>1020.7892216934413,
784=>1019.715761123694,
785=>1018.6416655766976,
786=>1017.5669375811376,
787=>1016.4915796671878,
788=>1015.415594366505,
789=>1014.338984212224,
790=>1013.261751738949,
791=>1012.1838994827508,
792=>1011.1054299811587,
793=>1010.0263457731553,
794=>1008.94664939917,
795=>1007.8663434010738,
796=>1006.7854303221728,
797=>1005.7039127072021,
798=>1004.6217931023203,
799=>1003.5390740551034,
800=>1002.455758114538,
801=>1001.3718478310163,
802=>1000.2873457563301,
803=>999.2022544436638,
804=>998.1165764475893,
805=>997.0303143240598,
806=>995.9434706304035,
807=>994.8560479253175,
808=>993.7680487688626,
809=>992.6794757224566,
810=>991.5903313488681,
811=>990.5006182122107,
812=>989.4103388779373,
813=>988.3194959128339,
814=>987.2280918850129,
815=>986.1361293639077,
816=>985.0436109202669,
817=>983.9505391261479,
818=>982.8569165549102,
819=>981.7627457812106,
820=>980.6680293809961,
821=>979.5727699314984,
822=>978.4769700112279,
823=>977.3806321999668,
824=>976.2837590787642,
825=>975.1863532299292,
826=>974.0884172370254,
827=>972.9899536848637,
828=>971.8909651594979,
829=>970.7914542482172,
830=>969.6914235395407,
831=>968.5908756232113,
832=>967.4898130901897,
833=>966.3882385326476,
834=>965.2861545439629,
835=>964.183563718712,
836=>963.0804686526653,
837=>961.9768719427798,
838=>960.8727761871934,
839=>959.7681839852196,
840=>958.6630979373396,
841=>957.5575206451981,
842=>956.451454711596,
843=>955.3449027404846,
844=>954.2378673369593,
845=>953.1303511072539,
846=>952.022356658734,
847=>950.9138865998912,
848=>949.8049435403364,
849=>948.6955300907945,
850=>947.5856488630977,
851=>946.4753024701795,
852=>945.3644935260685,
853=>944.2532246458819,
854=>943.1414984458202,
855=>942.0293175431605,
856=>940.9166845562497,
857=>939.8036021045001,
858=>938.6900728083815,
859=>937.5760992894154,
860=>936.46168417017,
861=>935.3468300742522,
862=>934.2315396263032,
863=>933.1158154519906,
864=>931.9996601780039,
865=>930.8830764320472,
866=>929.7660668428331,
867=>928.6486340400769,
868=>927.5307806544906,
869=>926.4125093177759,
870=>925.2938226626184,
871=>924.1747233226819,
872=>923.0552139326016,
873=>921.935297127978,
874=>920.8149755453703,
875=>919.6942518222918,
876=>918.573128597201,
877=>917.4516085094986,
878=>916.3296941995181,
879=>915.2073883085224,
880=>914.0846934786948,
881=>912.9616123531359,
882=>911.8381475758546,
883=>910.7143017917633,
884=>909.5900776466715,
885=>908.4654777872796,
886=>907.3405048611719,
887=>906.2151615168116,
888=>905.0894504035339,
889=>903.9633741715394,
890=>902.8369354718886,
891=>901.7101369564956,
892=>900.5829812781209,
893=>899.4554710903664,
894=>898.3276090476684,
895=>897.1993978052917,
896=>896.070840019323,
897=>894.941938346665,
898=>893.8126954450299,
899=>892.6831139729331,
900=>891.5531965896876,
901=>890.4229459553967,
902=>889.2923647309482,
903=>888.1614555780087,
904=>887.0302211590165,
905=>885.8986641371757,
906=>884.7667871764497,
907=>883.6345929415555,
908=>882.502084097957,
909=>881.369263311858,
910=>880.2361332501978,
911=>879.1026965806433,
912=>877.968955971583,
913=>876.834914092121,
914=>875.7005736120716,
915=>874.5659372019506,
916=>873.4310075329714,
917=>872.295787277038,
918=>871.1602791067377,
919=>870.024485695336,
920=>868.8884097167704,
921=>867.752053845643,
922=>866.6154207572149,
923=>865.4785131274002,
924=>864.3413336327591,
925=>863.2038849504918,
926=>862.0661697584322,
927=>860.9281907350421,
928=>859.7899505594037,
929=>858.6514519112143,
930=>857.51269747078,
931=>856.3736899190092,
932=>855.2344319374051,
933=>854.0949262080617,
934=>852.9551754136559,
935=>851.8151822374409,
936=>850.6749493632417,
937=>849.5344794754467,
938=>848.3937752590024,
939=>847.2528393994072,
940=>846.111674582705,
941=>844.9702834954784,
942=>843.8286688248426,
943=>842.6868332584395,
944=>841.5447794844308,
945=>840.4025101914923,
946=>839.2600280688066,
947=>838.1173358060579,
948=>836.9744360934246,
949=>835.831331621574,
950=>834.6880250816552,
951=>833.5445191652927,
952=>832.4008165645812,
953=>831.2569199720776,
954=>830.1128320807964,
955=>828.9685555842011,
956=>827.8240931762007,
957=>826.679447551141,
958=>825.5346214037994,
959=>824.3896174293782,
960=>823.2444383234987,
961=>822.0990867821937,
962=>820.9535655019029,
963=>819.807877179465,
964=>818.6620245121123,
965=>817.5160101974637,
966=>816.3698369335189,
967=>815.2235074186517,
968=>814.0770243516035,
969=>812.9303904314778,
970=>811.7836083577329,
971=>810.6366808301757,
972=>809.4896105489557,
973=>808.3424002145587,
974=>807.1950525278,
975=>806.0475701898183,
976=>804.8999559020691,
977=>803.752212366319,
978=>802.6043422846384,
979=>801.4563483593959,
980=>800.3082332932518,
981=>799.1599997891511,
982=>798.011650550318,
983=>796.8631882802493,
984=>795.7146156827074,
985=>794.5659354617148,
986=>793.4171503215475,
987=>792.2682629667281,
988=>791.11927610202,
989=>789.9701924324211,
990=>788.8210146631571,
991=>787.6717454996749,
992=>786.5223876476368,
993=>785.3729438129144,
994=>784.2234167015805,
995=>783.0738090199052,
996=>781.9241234743478,
997=>780.7743627715506,
998=>779.6245296183332,
999=>778.4746267216857,
1000=>777.3246567887627,
1001=>776.1746225268759,
1002=>775.0245266434888,
1003=>773.8743718462105,
1004=>772.7241608427878,
1005=>771.5738963411006,
1006=>770.4235810491544,
1007=>769.2732176750746,
1008=>768.1228089270992,
1009=>766.9723575135737,
1010=>765.8218661429435,
1011=>764.6713375237483,
1012=>763.5207743646157,
1013=>762.3701793742543,
1014=>761.2195552614477,
1015=>760.068904735048,
1016=>758.91823050397,
1017=>757.7675352771834,
1018=>756.6168217637079,
1019=>755.4660926726065,
1020=>754.3153507129782,
1021=>753.1645985939529,
1022=>752.0138390246839,
1023=>750.8630747143427,
1024=>749.7123083721111,
1025=>748.5615427071764,
1026=>747.4107804287241,
1027=>746.2600242459315,
1028=>745.1092768679619,
1029=>743.9585410039576,
1030=>742.8078193630339,
1031=>741.6571146542725,
1032=>740.5064295867156,
1033=>739.3557668693588,
1034=>738.2051292111452,
1035=>737.0545193209587,
1036=>735.9039399076183,
1037=>734.7533936798708,
1038=>733.602883346385,
1039=>732.4524116157455,
1040=>731.3019811964455,
1041=>730.1515947968812,
1042=>729.0012551253453,
1043=>727.8509648900205,
1044=>726.7007267989725,
1045=>725.5505435601451,
1046=>724.4004178813526,
1047=>723.2503524702736,
1048=>722.1003500344449,
1049=>720.9504132812555,
1050=>719.8005449179389,
1051=>718.6507476515683,
1052=>717.5010241890493,
1053=>716.351377237114,
1054=>715.2018095023137,
1055=>714.052323691014,
1056=>712.902922509387,
1057=>711.7536086634055,
1058=>710.6043848588381,
1059=>709.4552538012393,
1060=>708.3062181959467,
1061=>707.1572807480729,
1062=>706.008444162499,
1063=>704.8597111438689,
1064=>703.7110843965828,
1065=>702.5625666247909,
1066=>701.4141605323861,
1067=>700.265868822999,
1068=>699.1176941999909,
1069=>697.969639366447,
1070=>696.8217070251711,
1071=>695.6738998786783,
1072=>694.5262206291886,
1073=>693.3786719786217,
1074=>692.2312566285891,
1075=>691.083977280389,
1076=>689.9368366349992,
1077=>688.7898373930707,
1078=>687.6429822549222,
1079=>686.4962739205326,
1080=>685.3497150895355,
1081=>684.2033084612123,
1082=>683.0570567344864,
1083=>681.9109626079162,
1084=>680.7650287796891,
1085=>679.6192579476157,
1086=>678.4736528091216,
1087=>677.3282160612438,
1088=>676.182950400622,
1089=>675.037858523493,
1090=>673.892943125685,
1091=>672.7482069026103,
1092=>671.60365254926,
1093=>670.4592827601961,
1094=>669.3151002295468,
1095=>668.1711076509994,
1096=>667.0273077177935,
1097=>665.8837031227156,
1098=>664.7402965580926,
1099=>663.5970907157842,
1100=>662.4540882871786,
1101=>661.3112919631845,
1102=>660.1687044342259,
1103=>659.0263283902344,
1104=>657.8841665206445,
1105=>656.7422215143863,
1106=>655.600496059879,
1107=>654.4589928450253,
1108=>653.3177145572046,
1109=>652.1766638832667,
1110=>651.0358435095254,
1111=>649.8952561217527,
1112=>648.754904405172,
1113=>647.6147910444515,
1114=>646.4749187236985,
1115=>645.3352901264532,
1116=>644.1959079356811,
1117=>643.0567748337686,
1118=>641.9178935025152,
1119=>640.7792666231273,
1120=>639.640896876213,
1121=>638.5027869417747,
1122=>637.3649394992032,
1123=>636.227357227271,
1124=>635.0900428041272,
1125=>633.952998907289,
1126=>632.8162282136378,
1127=>631.6797333994116,
1128=>630.5435171401983,
1129=>629.4075821109309,
1130=>628.2719309858797,
1131=>627.1365664386467,
1132=>626.0014911421595,
1133=>624.8667077686646,
1134=>623.7322189897211,
1135=>622.5980274761946,
1136=>621.464135898251,
1137=>620.3305469253503,
1138=>619.1972632262392,
1139=>618.0642874689466,
1140=>616.9316223207763,
1141=>615.7992704483005,
1142=>614.6672345173539,
1143=>613.5355171930278,
1144=>612.4041211396633,
1145=>611.2730490208446,
1146=>610.142303499394,
1147=>609.0118872373646,
1148=>607.8818028960342,
1149=>606.7520531358994,
1150=>605.622640616669,
1151=>604.4935679972581,
1152=>603.364837935781,
1153=>602.2364530895463,
1154=>601.1084161150495,
1155=>599.9807296679668,
1156=>598.8533964031496,
1157=>597.726418974618,
1158=>596.5998000355537,
1159=>595.4735422382951,
1160=>594.3476482343299,
1161=>593.2221206742898,
1162=>592.0969622079433,
1163=>590.9721754841903,
1164=>589.8477631510556,
1165=>588.723727855682,
1166=>587.6000722443255,
1167=>586.4767989623476,
1168=>585.35391065421,
1169=>584.231409963468,
1170=>583.1092995327642,
1171=>581.987582003823,
1172=>580.8662600174429,
1173=>579.7453362134919,
1174=>578.6248132309005,
1175=>577.5046937076551,
1176=>576.3849802807929,
1177=>575.2656755863948,
1178=>574.1467822595789,
1179=>573.0283029344957,
1180=>571.9102402443208,
1181=>570.7925968212487,
1182=>569.6753752964868,
1183=>568.5585783002493,
1184=>567.4422084617515,
1185=>566.3262684092018,
1186=>565.2107607697986,
1187=>564.0956881697207,
1188=>562.9810532341235,
1189=>561.8668585871318,
1190=>560.7531068518336,
1191=>559.6398006502748,
1192=>558.5269426034519,
1193=>557.4145353313066,
1194=>556.3025814527191,
1195=>555.1910835855025,
1196=>554.0800443463963,
1197=>552.9694663510599,
1198=>551.859352214067,
1199=>550.7497045488999,
1200=>549.6405259679416,
1201=>548.5318190824717,
1202=>547.4235865026586,
1203=>546.3158308375549,
1204=>545.2085546950894,
1205=>544.1017606820628,
1206=>542.9954514041406,
1207=>541.8896294658466,
1208=>540.7842974705579,
1209=>539.679458020498,
1210=>538.5751137167306,
1211=>537.4712671591537,
1212=>536.3679209464939,
1213=>535.2650776762996,
1214=>534.162739944935,
1215=>533.0609103475742,
1216=>531.9595914781955,
1217=>530.8587859295741,
1218=>529.758496293277,
1219=>528.6587251596568,
1220=>527.5594751178455,
1221=>526.4607487557475,
1222=>525.3625486600356,
1223=>524.2648774161427,
1224=>523.1677376082567,
1225=>522.0711318193149,
1226=>520.9750626309971,
1227=>519.8795326237195,
1228=>518.7845443766294,
1229=>517.6901004675984,
1230=>516.596203473217,
1231=>515.5028559687873,
1232=>514.4100605283188,
1233=>513.3178197245205,
1234=>512.2261361287958,
1235=>511.1350123112368,
1236=>510.0444508406172,
1237=>508.95445428438677,
1238=>507.86502520866566,
1239=>506.77616617823804,
1240=>505.68787975654595,
1241=>504.60016850568303,
1242=>503.51303498638936,
1243=>502.4264817580447,
1244=>501.34051137866237,
1245=>500.255126404884,
1246=>499.1703293919729,
1247=>498.0861228938078,
1248=>497.00250946287747,
1249=>495.91949165027495,
1250=>494.8370720056902,
1251=>493.75525307740537,
1252=>492.67403741228867,
1253=>491.59342755578723,
1254=>490.5134260519227,
1255=>489.4340354432845,
1256=>488.3552582710233,
1257=>487.277097074846,
1258=>486.1995543930095,
1259=>485.1226327623141,
1260=>484.04633471809825,
1261=>482.97066279423234,
1262=>481.8956195231129,
1263=>480.82120743565594,
1264=>479.7474290612918,
1265=>478.67428692795926,
1266=>477.6017835620985,
1267=>476.52992148864644,
1268=>475.45870323103014,
1269=>474.38813131116063,
1270=>473.3182082494278,
1271=>472.24893656469357,
1272=>471.18031877428683,
1273=>470.1123573939963,
1274=>469.04505493806596,
1275=>467.97841391918854,
1276=>466.91243684849894,
1277=>465.84712623556976,
1278=>464.7824845884041,
1279=>463.71851441343046,
1280=>462.65521821549606,
1281=>461.5925984978619,
1282=>460.53065776219626,
1283=>459.46939850856864,
1284=>458.4088232354445,
1285=>457.34893443967906,
1286=>456.289734616511,
1287=>455.23122625955733,
1288=>454.1734118608072,
1289=>453.11629391061604,
1290=>452.05987489769916,
1291=>451.0041573091271,
1292=>449.94914363031876,
1293=>448.89483634503557,
1294=>447.8412379353765,
1295=>446.7883508817714,
1296=>445.7361776629752,
1297=>444.6847207560625,
1298=>443.63398263642165,
1299=>442.5839657777488,
1300=>441.5346726520415,
1301=>440.48610572959404,
1302=>439.43826747899124,
1303=>438.3911603671016,
1304=>437.34478685907317,
1305=>436.2991494183263,
1306=>435.254250506549,
1307=>434.2100925836902,
1308=>433.16667810795457,
1309=>432.1240095357964,
1310=>431.0820893219144,
1311=>430.04091991924435,
1312=>429.00050377895553,
1313=>427.9608433504431,
1314=>426.92194108132406,
1315=>425.8837994174296,
1316=>424.84642080280094,
1317=>423.8098076796818,
1318=>422.77396248851494,
1319=>421.7388876679346,
1320=>420.70458565476156,
1321=>419.67105888399726,
1322=>418.6383097888181,
1323=>417.60634080056906,
1324=>416.5751543487592,
1325=>415.5447528610552,
1326=>414.5151387632755,
1327=>413.48631447938493,
1328=>412.4582824314891,
1329=>411.4310450398286,
1330=>410.40460472277215,
1331=>409.3789638968133,
1332=>408.3541249765627,
1333=>407.33009037474324,
1334=>406.3068625021844,
1335=>405.28444376781624,
1336=>404.26283657866423,
1337=>403.2420433398425,
1338=>402.22206645454963,
1339=>401.20290832406215,
1340=>400.184571347729,
1341=>399.1670579229659,
1342=>398.15037044525013,
1343=>397.1345113081135,
1344=>396.1194829031384,
1345=>395.1052876199517,
1346=>394.09192784621837,
1347=>393.07940596763666,
1348=>392.0677243679321,
1349=>391.0568854288524,
1350=>390.0468915301604,
1351=>389.0377450496306,
1352=>388.0294483630419,
1353=>387.0220038441729,
1354=>386.0154138647957,
1355=>385.00968079467077,
1356=>384.00480700154145,
1357=>383.00079485112724,
1358=>381.99764670712,
1359=>380.9953649311773,
1360=>379.9939518829168,
1361=>378.9934099199114,
1362=>377.9937413976828,
1363=>376.994948669697,
1364=>375.99703408735724,
1365=>375.00000000000017,
1366=>374.00384875488925,
1367=>373.0085826972096,
1368=>372.0142041700622,
1369=>371.02071551445925,
1370=>370.0281190693167,
1371=>369.0364171714511,
1372=>368.04561215557254,
1373=>367.05570635427995,
1374=>366.0667020980549,
1375=>365.07860171525687,
1376=>364.09140753211716,
1377=>363.10512187273366,
1378=>362.11974705906545,
1379=>361.13528541092734,
1380=>360.15173924598406,
1381=>359.1691108797455,
1382=>358.1874026255602,
1383=>357.2066167946109,
1384=>356.2267556959089,
1385=>355.24782163628817,
1386=>354.26981692040033,
1387=>353.29274385070903,
1388=>352.316604727485,
1389=>351.3414018487992,
1390=>350.36713751051934,
1391=>349.39381400630344,
1392=>348.42143362759435,
1393=>347.4499986636148,
1394=>346.47951140136155,
1395=>345.5099741256007,
1396=>344.5413891188609,
1397=>343.5737586614298,
1398=>342.60708503134754,
1399=>341.64137050440155,
1400=>340.6766173541215,
1401=>339.71282785177385,
1402=>338.7500042663556,
1403=>337.78814886459065,
1404=>336.8272639109232,
1405=>335.8673516675127,
1406=>334.9084143942289,
1407=>333.9504543486458,
1408=>332.99347378603744,
1409=>332.03747495937085,
1410=>331.0824601193027,
1411=>330.1284315141729,
1412=>329.17539138999956,
1413=>328.22334199047333,
1414=>327.27228555695285,
1415=>326.3222243284591,
1416=>325.3731605416694,
1417=>324.42509643091375,
1418=>323.47803422816816,
1419=>322.53197616305,
1420=>321.5869244628128,
1421=>320.6428813523406,
1422=>319.69984905414344,
1423=>318.7578297883509,
1424=>317.8168257727081,
1425=>316.87683922257014,
1426=>315.93787235089644,
1427=>314.99992736824623,
1428=>314.0630064827728,
1429=>313.12711190021787,
1430=>312.1922458239078,
1431=>311.25841045474726,
1432=>310.3256079912145,
1433=>309.393840629356,
1434=>308.46311056278125,
1435=>307.533419982658,
1436=>306.6047710777063,
1437=>305.67716603419404,
1438=>304.75060703593186,
1439=>303.8250962642675,
1440=>302.9006358980811,
1441=>301.97722811377963,
1442=>301.05487508529217,
1443=>300.13357898406474,
1444=>299.2133419790548,
1445=>298.29416623672694,
1446=>297.3760539210467,
1447=>296.45900719347674,
1448=>295.54302821297,
1449=>294.62811913596664,
1450=>293.71428211638766,
1451=>292.8015193056302,
1452=>291.88983285256245,
1453=>290.9792249035186,
1454=>290.069697602294,
1455=>289.16125309013927,
1456=>288.2538935057563,
1457=>287.34762098529285,
1458=>286.44243766233745,
1459=>285.53834566791414,
1460=>284.63534713047824,
1461=>283.7334441759099,
1462=>282.8326389275108,
1463=>281.93293350599805,
1464=>281.0343300294996,
1465=>280.136830613549,
1466=>279.2404373710807,
1467=>278.34515241242514,
1468=>277.4509778453028,
1469=>276.5579157748209,
1470=>275.66596830346714,
1471=>274.7751375311053,
1472=>273.8854255549702,
1473=>272.9968344696628,
1474=>272.1093663671451,
1475=>271.223023336735,
1476=>270.3378074651022,
1477=>269.4537208362627,
1478=>268.5707655315737,
1479=>267.6889436297294,
1480=>266.80825720675546,
1481=>265.92870833600443,
1482=>265.0502990881504,
1483=>264.1730315311849,
1484=>263.2969077304118,
1485=>262.4219297484418,
1486=>261.5480996451885,
1487=>260.67541947786304,
1488=>259.80389130096876,
1489=>258.9335171662975,
1490=>258.0642991229243,
1491=>257.19623921720205,
1492=>256.32933949275736,
1493=>255.46360199048553,
1494=>254.59902874854578,
1495=>253.73562180235564,
1496=>252.87338318458774,
1497=>252.01231492516393,
1498=>251.15241905125072,
1499=>250.29369758725448,
1500=>249.43615255481672,
1501=>248.57978597280976,
1502=>247.7245998573306,
1503=>246.870596221698,
1504=>246.01777707644635,
1505=>245.16614442932223,
1506=>244.3157002852783,
1507=>243.46644664646885,
1508=>242.61838551224605,
1509=>241.77151887915454,
1510=>240.92584874092654,
1511=>240.08137708847772,
1512=>239.23810590990206,
1513=>238.39603719046744,
1514=>237.55517291261037,
1515=>236.71551505593254,
1516=>235.87706559719504,
1517=>235.03982651031413,
1518=>234.2037997663565,
1519=>233.36898733353507,
1520=>232.53539117720322,
1521=>231.70301325985156,
1522=>230.8718555411025,
1523=>230.04191997770556,
1524=>229.21320852353347,
1525=>228.38572312957683,
1526=>227.55946574393988,
1527=>226.73443831183545,
1528=>225.9106427755812,
1529=>225.08808107459447,
1530=>224.26675514538795,
1531=>223.44666692156477,
1532=>222.6278183338144,
1533=>221.81021130990814,
1534=>220.99384777469345,
1535=>220.1787296500912,
1536=>219.36485885509012,
1537=>218.5522373057421,
1538=>217.7408669151581,
1539=>216.93074959350395,
1540=>216.12188724799466,
1541=>215.31428178289138,
1542=>214.50793509949597,
1543=>213.70284909614702,
1544=>212.8990256682149,
1545=>212.09646670809764,
1546=>211.2951741052168,
1547=>210.49514974601175,
1548=>209.69639551393698,
1549=>208.89891328945635,
1550=>208.10270495003908,
1551=>207.3077723701556,
1552=>206.51411742127277,
1553=>205.72174197184972,
1554=>204.93064788733273,
1555=>204.14083703015217,
1556=>203.352311259717,
1557=>202.56507243241083,
1558=>201.77912240158764,
1559=>200.994463017567,
1560=>200.2110961276304,
1561=>199.42902357601588,
1562=>198.6482472039146,
1563=>197.86876884946628,
1564=>197.09059034775476,
1565=>196.31371353080374,
1566=>195.5381402275724,
1567=>194.7638722639507,
1568=>193.99091146275612,
1569=>193.21925964372838,
1570=>192.44891862352597,
1571=>191.67989021572112,
1572=>190.9121762307958,
1573=>190.14577847613737,
1574=>189.3806987560348,
1575=>188.61693887167405,
1576=>187.85450062113387,
1577=>187.09338579938105,
1578=>186.33359619826763,
1579=>185.57513360652467,
1580=>184.81799980976018,
1581=>184.06219659045303,
1582=>183.3077257279499,
1583=>182.5545889984611,
1584=>181.8027881750554,
1585=>181.0523250276575,
1586=>180.30320132304155,
1587=>179.5554188248292,
1588=>178.8089792934844,
1589=>178.0638844863097,
1590=>177.3201361574413,
1591=>176.57773605784587,
1592=>175.83668593531593,
1593=>175.09698753446537,
1594=>174.35864259672644,
1595=>173.62165286034485,
1596=>172.88602006037547,
1597=>172.15174592867913,
1598=>171.41883219391786,
1599=>170.68728058155045,
1600=>169.9570928138296,
1601=>169.22827060979682,
1602=>168.50081568527912,
1603=>167.774729752884,
1604=>167.05001452199656,
1605=>166.32667169877493,
1606=>165.60470298614564,
1607=>164.8841100838007,
1608=>164.16489468819327,
1609=>163.4470584925332,
1610=>162.73060318678336,
1611=>162.01553045765593,
1612=>161.30184198860832,
1613=>160.58953945983808,
1614=>159.87862454828098,
1615=>159.16909892760555,
1616=>158.46096426820952,
1617=>157.75422223721625,
1618=>157.04887449847035,
1619=>156.34492271253384,
1620=>155.64236853668228,
1621=>154.94121362490114,
1622=>154.24145962788145,
1623=>153.54310819301634,
1624=>152.84616096439686,
1625=>152.15061958280842,
1626=>151.45648568572608,
1627=>150.76376090731208,
1628=>150.07244687841091,
1629=>149.38254522654586,
1630=>148.69405757591505,
1631=>148.0069855473879,
1632=>147.32133075850095,
1633=>146.63709482345416,
1634=>145.95427935310727,
1635=>145.2728859549759,
1636=>144.5929162332277,
1637=>143.91437178867886,
1638=>143.23725421878953,
1639=>142.5615651176612,
1640=>141.88730607603213,
1641=>141.21447868127427,
1642=>140.54308451738848,
1643=>139.87312516500197,
1644=>139.20460220136408,
1645=>138.53751720034177,
1646=>137.8718717324175,
1647=>137.20766736468454,
1648=>136.54490566084314,
1649=>135.88358818119764,
1650=>135.22371648265187,
1651=>134.56529211870645,
1652=>133.9083166394538,
1653=>133.25279159157606,
1654=>132.59871851834043,
1655=>131.94609895959582,
1656=>131.29493445176934,
1657=>130.6452265278624,
1658=>129.99697671744696,
1659=>129.3501865466627,
1660=>128.70485753821288,
1661=>128.06099121136083,
1662=>127.41858908192592,
1663=>126.77765266228107,
1664=>126.13818346134849,
1665=>125.50018298459531,
1666=>124.86365273403203,
1667=>124.22859420820748,
1668=>123.59500890220545,
1669=>122.9628983076417,
1670=>122.3322639126601,
1671=>121.70310720192936,
1672=>121.07542965663868,
1673=>120.4492327544956,
1674=>119.82451796972168,
1675=>119.20128677304922,
1676=>118.57954063171769,
1677=>117.9592810094706,
1678=>117.34050936655171,
1679=>116.72322715970142,
1680=>116.10743584215402,
1681=>115.49313686363371,
1682=>114.88033167035144,
1683=>114.26902170500148,
1684=>113.65920840675778,
1685=>113.05089321127082,
1686=>112.44407755066413,
1687=>111.8387628535313,
1688=>111.23495054493173,
1689=>110.63264204638824,
1690=>110.03183877588333,
1691=>109.43254214785566,
1692=>108.83475357319674,
1693=>108.23847445924798,
1694=>107.64370620979707,
1695=>107.05045022507488,
1696=>106.45870790175206,
1697=>105.86848063293519,
1698=>105.27976980816482,
1699=>104.69257681341094,
1700=>104.10690303107026,
1701=>103.52274983996301,
1702=>102.94011861532942,
1703=>102.35901072882689,
1704=>101.77942754852597,
1705=>101.20137043890838,
1706=>100.62484076086253,
1707=>100.04983987168123,
1708=>99.476369125058,
1709=>98.90442987108406,
1710=>98.33402345624518,
1711=>97.76515122341812,
1712=>97.19781451186816,
1713=>96.63201465724558,
1714=>96.06775299158232,
1715=>95.50503084328932,
1716=>94.9438495371528,
1717=>94.38421039433149,
1718=>93.82611473235374,
1719=>93.26956386511392,
1720=>92.71455910286977,
1721=>92.16110175223912,
1722=>91.60919311619648,
1723=>91.058834494071,
1724=>90.51002718154166,
1725=>89.96277247063608,
1726=>89.41707164972672,
1727=>88.87292600352714,
1728=>88.33033681309041,
1729=>87.7893053558048,
1730=>87.2498329053916,
1731=>86.71192073190127,
1732=>86.17557010171174,
1733=>85.6407822775243,
1734=>85.10755851836086,
1735=>84.5759000795615,
1736=>84.04580821278103,
1737=>83.51728416598576,
1738=>82.99032918345165,
1739=>82.46494450576006,
1740=>81.94113136979604,
1741=>81.41889100874437,
1742=>80.89822465208749,
1743=>80.37913352560201,
1744=>79.86161885135607,
1745=>79.3456818477066,
1746=>78.83132372929606,
1747=>78.31854570705025,
1748=>77.80734898817457,
1749=>77.29773477615186,
1750=>76.78970427073966,
1751=>76.28325866796615,
1752=>75.77839916012931,
1753=>75.27512693579251,
1754=>74.77344317978225,
1755=>74.27334907318573,
1756=>73.77484579334725,
1757=>73.2779345138664,
1758=>72.78261640459436,
1759=>72.28889263163182,
1760=>71.79676435732597,
1761=>71.306232740268,
1762=>70.81729893529007,
1763=>70.32996409346231,
1764=>69.84422936209091,
1765=>69.36009588471507,
1766=>68.87756480110386,
1767=>68.39663724725449,
1768=>67.91731435538838,
1769=>67.43959725394984,
1770=>66.96348706760216,
1771=>66.48898491722593,
1772=>66.01609191991588,
1773=>65.54480918897855,
1774=>65.07513783392938,
1775=>64.60707896049053,
1776=>64.14063367058725,
1777=>63.67580306234663,
1778=>63.212588230094525,
1779=>62.75099026435237,
1780=>62.29101025183536,
1781=>61.832649275449626,
1782=>61.375908414289825,
1783=>60.92078874363585,
1784=>60.467291334951824,
1785=>60.01541725588186,
1786=>59.56516757024883,
1787=>59.11654333805143,
1788=>58.66954561546129,
1789=>58.22417545482108,
1790=>57.78043390464143,
1791=>57.33832200959944,
1792=>56.89784081053506,
1793=>56.4589913444496,
1794=>56.02177464450244,
1795=>55.58619174000955,
1796=>55.15224365643985,
1797=>54.71993141541395,
1798=>54.28925603470145,
1799=>53.860218528217956,
1800=>53.43281990602327,
1801=>53.007061174319006,
1802=>52.582943335445975,
1803=>52.16046738788168,
1804=>51.73963432623873,
1805=>51.3204451412613,
1806=>50.902900819824254,
1807=>50.48700234492924,
1808=>50.07275069570392,
1809=>49.66014684739855,
1810=>49.24919177138372,
1811=>48.83988643514908,
1812=>48.43223180229995,
1813=>48.02622883255583,
1814=>47.62187848174733,
1815=>47.219181701814705,
1816=>46.81813944080557,
1817=>46.41875264287148,
1818=>46.0210222482674,
1819=>45.6249491933487,
1820=>45.230534410568794,
1821=>44.83777882847687,
1822=>44.446683371716404,
1823=>44.05724896102208,
1824=>43.669476513218456,
1825=>43.283366941217196,
1826=>42.89892115401517,
1827=>42.51614005669262,
1828=>42.13502455041021,
1829=>41.75557553240742,
1830=>41.37779389600075,
1831=>41.00168053058121,
1832=>40.62723632161192,
1833=>40.254462150626864,
1834=>39.88335889522807,
1835=>39.51392742908388,
1836=>39.146168621926904,
1837=>38.78008333955165,
1838=>38.41567244381315,
1839=>38.05293679262422,
1840=>37.69187723995378,
1841=>37.3324946358249,
1842=>36.97478982631253,
1843=>36.61876365354192,
1844=>36.26441695568599,
1845=>35.91175056696443,
1846=>35.56076531764029,
1847=>35.21146203401952,
1848=>34.86384153844779,
1849=>34.517904649309344,
1850=>34.17365218102452,
1851=>33.83108494404837,
1852=>33.49020374486861,
1853=>33.15100938600335,
1854=>32.81350266599975,
1855=>32.47768437943114,
1856=>32.14355531689682,
1857=>31.81111626501854,
1858=>31.48036800643979,
1859=>31.151311319823208,
1860=>30.823946979849325,
1861=>30.498275757214287,
1862=>30.17429841862804,
1863=>29.85201572681308,
1864=>29.53142844050228,
1865=>29.21253731443676,
1866=>28.895343099364823,
1867=>28.579846542039604,
1868=>28.266048385217687,
1869=>27.953949367656946,
1870=>27.64355022411553,
1871=>27.334851685349122,
1872=>27.027854478110044,
1873=>26.722559325145312,
1874=>26.41896694519494,
1875=>26.117078052989882,
1876=>25.816893359250912,
1877=>25.518413570686448,
1878=>25.22163938999165,
1879=>24.92657151584592,
1880=>24.633210642911422,
1881=>24.341557461832053,
1882=>24.051612659230727,
1883=>23.76337691770925,
1884=>23.476850915845375,
1885=>23.19203532819165,
1886=>22.90893082527407,
1887=>22.627538073590358,
1888=>22.347857735608272,
1889=>22.069890469764005,
1890=>21.793636930460934,
1891=>21.519097768067923,
1892=>21.24627362891772,
1893=>20.975165155305376,
1894=>20.705772985486874,
1895=>20.438097753677766,
1896=>20.17214009005113,
1897=>19.907900620737223,
1898=>19.645379967820304,
1899=>19.384578749338743,
1900=>19.125497579282865,
1901=>18.86813706759324,
1902=>18.61249782016,
1903=>18.358580438820695,
1904=>18.106385521359357,
1905=>17.85591366150493,
1906=>17.607165448929663,
1907=>17.36014146924822,
1908=>17.11484230401561,
1909=>16.871268530726525,
1910=>16.629420722813506,
1911=>16.389299449645705,
1912=>16.15090527652785,
1913=>15.914238764698439,
1914=>15.679300471328474,
1915=>15.44609094952068,
1916=>15.21461074830745,
1917=>14.984860412650278,
1918=>14.75684048343794,
1919=>14.530551497485476,
1920=>14.305993987532815,
1921=>14.083168482243423,
1922=>13.862075506203496,
1923=>13.64271557992015,
1924=>13.425089219820848,
1925=>13.209196938251466,
1926=>12.99503924347539,
1927=>12.78261663967271,
1928=>12.571929626938527,
1929=>12.362978701281577,
1930=>12.155764354624012,
1931=>11.950287074799462,
1932=>11.746547345551676,
1933=>11.544545646534402,
1934=>11.34428245330912,
1935=>11.145758237344694,
1936=>10.948973466016014,
1937=>10.753928602602741,
1938=>10.560624106288628,
1939=>10.369060432159927,
1940=>10.17923803120459,
1941=>9.991157350311369,
1942=>9.80481883226821,
1943=>9.620222915762042,
1944=>9.437370035377171,
1945=>9.256260621593924,
1946=>9.076895100788647,
1947=>8.899273895231886,
1948=>8.723397423087476,
1949=>8.54926609841209,
1950=>8.376880331153643,
1951=>8.206240527150499,
1952=>8.037347088131014,
1953=>7.870200411711608,
1954=>7.7048008913968715,
1955=>7.541148916577981,
1956=>7.379244872531672,
1957=>7.219089140420124,
1958=>7.060682097289373,
1959=>6.904024116068399,
1960=>6.7491155655686725,
1961=>6.595956810483017,
1962=>6.444548211384927,
1963=>6.294890124727317,
1964=>6.146982902842296,
1965=>6.0008268939396885,
1966=>5.856422442106918,
1967=>5.713769887307308,
1968=>5.5728695653803015,
1969=>5.433721808039877,
1970=>5.296326942873975,
1971=>5.160685293343931,
1972=>5.026797178783568,
1973=>4.894662914398509,
1974=>4.764282811265275,
1975=>4.63565717633071,
1976=>4.508786312411075,
1977=>4.3836705181918205,
1978=>4.260310088225992,
1979=>4.138705312934803,
1980=>4.018856478605585,
1981=>3.900763867391788,
1982=>3.7844277573127556,
1983=>3.66984842225213,
1984=>3.5570261319579686,
1985=>3.4459611520417184,
1986=>3.3366537439776494,
1987=>3.2291041651020578,
1988=>3.12331266861338,
1989=>3.019279503570715,
1990=>2.9170049148938233,
1991=>2.8164891433619914,
1992=>2.717732425614372,
1993=>2.6207349941485063,
1994=>2.525497077319983,
1995=>2.4320188993425518,
1996=>2.3403006802866457,
1997=>2.250342636079722,
1998=>2.162144978504898,
1999=>2.0757079152014057,
2000=>1.991031649663114,
2001=>1.9081163812389832,
2002=>1.826962305131815,
2003=>1.7475696123983653,
2004=>1.6699384899484357,
2005=>1.5940691205449866,
2006=>1.5199616828030003,
2007=>1.4476163511897084,
2008=>1.3770332960236829,
2009=>1.3082126834749488,
2010=>1.2411546755640757,
2011=>1.1758594301622907,
2012=>1.112327100990342,
2013=>1.0505578376191806,
2014=>0.9905517854688242,
2015=>0.9323090858082423,
2016=>0.8758298757550165,
2017=>0.8211142882752256,
2018=>0.7681624521827644,
2019=>0.7169744921393431,
2020=>0.6675505286539192,
2021=>0.6198906780826974,
2022=>0.5739950526285611,
2023=>0.5298637603414136,
2024=>0.48749690511692734,
2025=>0.44689458669722626,
2026=>0.40805690066986244,
2027=>0.37098393846883937,
2028=>0.33567578737245185,
2029=>0.302132530505105,
2030=>0.2703542468359501,
2031=>0.24034101117865703,
2032=>0.21209289419186916,
2033=>0.18560996237852123,
2034=>0.16089227808618034,
2035=>0.1379398995060228,
2036=>0.11675288067374368,
2037=>0.09733127146898823,
2038=>0.07967511761466994,
2039=>0.06378446067799359,
2040=>0.04965933806931844,
2041=>0.03729978304272663,
2042=>0.02670582469556848,
2043=>0.017877487968803507,
2044=>0.010814793646204635,
2045=>0.005517758355381375,
2046=>0.001986394566756644,
2047=>0.0002207105940215115,
2048=>0.0002207105940215115,
2049=>0.001986394566756644,
2050=>0.005517758355381375,
2051=>0.010814793646204635,
2052=>0.017877487968803507,
2053=>0.02670582469556848,
2054=>0.03729978304272663,
2055=>0.04965933806931844,
2056=>0.06378446067799359,
2057=>0.07967511761466994,
2058=>0.09733127146898823,
2059=>0.11675288067374368,
2060=>0.1379398995060228,
2061=>0.16089227808618034,
2062=>0.18560996237852123,
2063=>0.21209289419186916,
2064=>0.24034101117865703,
2065=>0.2703542468358364,
2066=>0.302132530505105,
2067=>0.33567578737245185,
2068=>0.3709839384687257,
2069=>0.40805690066986244,
2070=>0.44689458669722626,
2071=>0.48749690511692734,
2072=>0.5298637603414136,
2073=>0.5739950526285611,
2074=>0.6198906780826974,
2075=>0.6675505286539192,
2076=>0.7169744921393431,
2077=>0.7681624521827644,
2078=>0.8211142882752256,
2079=>0.8758298757550165,
2080=>0.9323090858082423,
2081=>0.9905517854688242,
2082=>1.0505578376191806,
2083=>1.112327100990342,
2084=>1.1758594301622907,
2085=>1.2411546755640757,
2086=>1.3082126834749488,
2087=>1.3770332960236829,
2088=>1.4476163511897084,
2089=>1.5199616828030003,
2090=>1.5940691205449866,
2091=>1.6699384899484357,
2092=>1.7475696123982516,
2093=>1.826962305131815,
2094=>1.9081163812389832,
2095=>1.991031649663114,
2096=>2.075707915201292,
2097=>2.162144978504898,
2098=>2.2503426360796084,
2099=>2.3403006802866457,
2100=>2.432018899342438,
2101=>2.525497077319983,
2102=>2.6207349941483926,
2103=>2.717732425614372,
2104=>2.8164891433619914,
2105=>2.9170049148937096,
2106=>3.019279503570715,
2107=>3.12331266861338,
2108=>3.229104165101944,
2109=>3.3366537439775357,
2110=>3.4459611520417184,
2111=>3.5570261319579686,
2112=>3.66984842225213,
2113=>3.7844277573127556,
2114=>3.900763867391788,
2115=>4.018856478605585,
2116=>4.138705312934803,
2117=>4.260310088226106,
2118=>4.3836705181918205,
2119=>4.508786312411075,
2120=>4.63565717633071,
2121=>4.764282811265275,
2122=>4.894662914398509,
2123=>5.026797178783568,
2124=>5.160685293343931,
2125=>5.296326942873975,
2126=>5.433721808039877,
2127=>5.572869565380415,
2128=>5.713769887307421,
2129=>5.856422442106918,
2130=>6.0008268939396885,
2131=>6.146982902842296,
2132=>6.294890124727317,
2133=>6.444548211384927,
2134=>6.5959568104831305,
2135=>6.7491155655686725,
2136=>6.904024116068399,
2137=>7.060682097289373,
2138=>7.219089140420124,
2139=>7.379244872531785,
2140=>7.541148916577981,
2141=>7.704800891396985,
2142=>7.870200411711608,
2143=>8.037347088131014,
2144=>8.206240527150499,
2145=>8.376880331153643,
2146=>8.54926609841209,
2147=>8.723397423087476,
2148=>8.899273895231772,
2149=>9.076895100788647,
2150=>9.256260621593924,
2151=>9.437370035377057,
2152=>9.620222915762042,
2153=>9.80481883226821,
2154=>9.991157350311255,
2155=>10.17923803120459,
2156=>10.369060432159927,
2157=>10.560624106288515,
2158=>10.753928602602741,
2159=>10.948973466016014,
2160=>11.145758237344694,
2161=>11.34428245330912,
2162=>11.544545646534289,
2163=>11.746547345551676,
2164=>11.950287074799348,
2165=>12.155764354624012,
2166=>12.362978701281577,
2167=>12.571929626938413,
2168=>12.78261663967271,
2169=>12.99503924347539,
2170=>13.209196938251353,
2171=>13.425089219820848,
2172=>13.64271557992015,
2173=>13.862075506203496,
2174=>14.083168482243423,
2175=>14.305993987532702,
2176=>14.530551497485476,
2177=>14.75684048343794,
2178=>14.984860412650278,
2179=>15.21461074830745,
2180=>15.44609094952068,
2181=>15.679300471328474,
2182=>15.914238764698439,
2183=>16.15090527652785,
2184=>16.389299449645705,
2185=>16.629420722813506,
2186=>16.871268530726525,
2187=>17.11484230401561,
2188=>17.36014146924822,
2189=>17.607165448929663,
2190=>17.855913661504815,
2191=>18.106385521359357,
2192=>18.35858043882058,
2193=>18.612497820159888,
2194=>18.868137067593125,
2195=>19.12549757928275,
2196=>19.38457874933863,
2197=>19.645379967820304,
2198=>19.90790062073711,
2199=>20.17214009005113,
2200=>20.438097753677653,
2201=>20.70577298548676,
2202=>20.975165155305262,
2203=>21.246273628917606,
2204=>21.519097768067923,
2205=>21.793636930460934,
2206=>22.06989046976389,
2207=>22.34785773560816,
2208=>22.627538073590358,
2209=>22.908930825273956,
2210=>23.192035328191423,
2211=>23.476850915845148,
2212=>23.763376917709138,
2213=>24.051612659230614,
2214=>24.341557461831826,
2215=>24.63321064291131,
2216=>24.926571515845808,
2217=>25.22163938999165,
2218=>25.518413570686448,
2219=>25.816893359250685,
2220=>26.11707805298977,
2221=>26.418966945194825,
2222=>26.722559325145312,
2223=>27.02785447810993,
2224=>27.334851685348895,
2225=>27.643550224115415,
2226=>27.953949367656946,
2227=>28.266048385217573,
2228=>28.57984654203949,
2229=>28.895343099364823,
2230=>29.212537314436645,
2231=>29.531428440502054,
2232=>29.852015726812965,
2233=>30.174298418627814,
2234=>30.49827575721406,
2235=>30.82394697984921,
2236=>31.151311319823094,
2237=>31.480368006439676,
2238=>31.811116265018427,
2239=>32.143555316896595,
2240=>32.477684379431025,
2241=>32.813502665999636,
2242=>33.151009386003466,
2243=>33.49020374486872,
2244=>33.831084944048484,
2245=>34.17365218102452,
2246=>34.517904649309344,
2247=>34.86384153844779,
2248=>35.21146203401952,
2249=>35.5607653176404,
2250=>35.91175056696443,
2251=>36.2644169556861,
2252=>36.61876365354192,
2253=>36.97478982631253,
2254=>37.33249463582479,
2255=>37.69187723995378,
2256=>38.05293679262422,
2257=>38.41567244381315,
2258=>38.78008333955165,
2259=>39.146168621926904,
2260=>39.51392742908388,
2261=>39.88335889522796,
2262=>40.254462150626864,
2263=>40.62723632161192,
2264=>41.00168053058121,
2265=>41.37779389600087,
2266=>41.75557553240753,
2267=>42.135024550410094,
2268=>42.51614005669262,
2269=>42.898921154015284,
2270=>43.28336694121731,
2271=>43.669476513218456,
2272=>44.05724896102208,
2273=>44.44668337171629,
2274=>44.83777882847676,
2275=>45.23053441056868,
2276=>45.6249491933487,
2277=>46.0210222482674,
2278=>46.41875264287137,
2279=>46.81813944080545,
2280=>47.219181701814705,
2281=>47.62187848174733,
2282=>48.02622883255572,
2283=>48.43223180229995,
2284=>48.83988643514908,
2285=>49.24919177138361,
2286=>49.66014684739844,
2287=>50.0727506957038,
2288=>50.48700234492924,
2289=>50.90290081982414,
2290=>51.32044514126119,
2291=>51.739634326238615,
2292=>52.16046738788168,
2293=>52.582943335445975,
2294=>53.00706117431889,
2295=>53.432819906023155,
2296=>53.86021852821784,
2297=>54.28925603470134,
2298=>54.71993141541395,
2299=>55.15224365643974,
2300=>55.58619174000944,
2301=>56.02177464450244,
2302=>56.45899134444949,
2303=>56.89784081053506,
2304=>57.338322009599324,
2305=>57.78043390464143,
2306=>58.224175454820966,
2307=>58.669545615461175,
2308=>59.116543338051315,
2309=>59.56516757024883,
2310=>60.01541725588186,
2311=>60.46729133495171,
2312=>60.92078874363585,
2313=>61.37590841428971,
2314=>61.832649275449626,
2315=>62.291010251835246,
2316=>62.750990264352254,
2317=>63.21258823009441,
2318=>63.67580306234663,
2319=>64.14063367058714,
2320=>64.60707896049041,
2321=>65.07513783392938,
2322=>65.54480918897855,
2323=>66.01609191991577,
2324=>66.48898491722582,
2325=>66.96348706760216,
2326=>67.43959725394984,
2327=>67.91731435538838,
2328=>68.39663724725438,
2329=>68.87756480110386,
2330=>69.36009588471495,
2331=>69.84422936209091,
2332=>70.3299640934622,
2333=>70.81729893528995,
2334=>71.30623274026789,
2335=>71.79676435732586,
2336=>72.2888926316316,
2337=>72.78261640459414,
2338=>73.27793451386617,
2339=>73.77484579334714,
2340=>74.27334907318561,
2341=>74.77344317978213,
2342=>75.27512693579229,
2343=>75.77839916012908,
2344=>76.28325866796604,
2345=>76.78970427073943,
2346=>77.29773477615186,
2347=>77.80734898817445,
2348=>78.31854570705002,
2349=>78.83132372929583,
2350=>79.34568184770637,
2351=>79.86161885135584,
2352=>80.3791335256019,
2353=>80.89822465208738,
2354=>81.41889100874414,
2355=>81.9411313697957,
2356=>82.46494450575983,
2357=>82.99032918345142,
2358=>83.51728416598553,
2359=>84.04580821278068,
2360=>84.57590007956139,
2361=>85.10755851836063,
2362=>85.64078227752395,
2363=>86.17557010171151,
2364=>86.71192073190105,
2365=>87.24983290539137,
2366=>87.78930535580469,
2367=>88.3303368130903,
2368=>88.87292600352691,
2369=>89.41707164972672,
2370=>89.9627724706362,
2371=>90.51002718154166,
2372=>91.05883449407088,
2373=>91.6091931161966,
2374=>92.16110175223923,
2375=>92.71455910286988,
2376=>93.26956386511404,
2377=>93.82611473235386,
2378=>94.38421039433138,
2379=>94.94384953715269,
2380=>95.50503084328932,
2381=>96.06775299158244,
2382=>96.63201465724569,
2383=>97.19781451186827,
2384=>97.76515122341823,
2385=>98.33402345624506,
2386=>98.90442987108418,
2387=>99.47636912505811,
2388=>100.04983987168134,
2389=>100.62484076086264,
2390=>101.2013704389085,
2391=>101.77942754852609,
2392=>102.35901072882677,
2393=>102.94011861532942,
2394=>103.52274983996313,
2395=>104.10690303107037,
2396=>104.69257681341105,
2397=>105.27976980816493,
2398=>105.86848063293519,
2399=>106.45870790175195,
2400=>107.05045022507488,
2401=>107.64370620979707,
2402=>108.23847445924787,
2403=>108.83475357319662,
2404=>109.43254214785554,
2405=>110.03183877588322,
2406=>110.63264204638813,
2407=>111.23495054493162,
2408=>111.8387628535312,
2409=>112.44407755066402,
2410=>113.0508932112707,
2411=>113.65920840675778,
2412=>114.26902170500136,
2413=>114.88033167035144,
2414=>115.4931368636336,
2415=>116.1074358421539,
2416=>116.72322715970131,
2417=>117.34050936655171,
2418=>117.95928100947049,
2419=>118.57954063171758,
2420=>119.2012867730491,
2421=>119.82451796972157,
2422=>120.44923275449548,
2423=>121.07542965663856,
2424=>121.70310720192924,
2425=>122.3322639126601,
2426=>122.9628983076417,
2427=>123.59500890220545,
2428=>124.22859420820737,
2429=>124.86365273403192,
2430=>125.5001829845952,
2431=>126.13818346134826,
2432=>126.77765266228107,
2433=>127.4185890819258,
2434=>128.06099121136072,
2435=>128.70485753821276,
2436=>129.3501865466626,
2437=>129.99697671744673,
2438=>130.64522652786218,
2439=>131.2949344517691,
2440=>131.9460989595957,
2441=>132.59871851834032,
2442=>133.25279159157594,
2443=>133.9083166394537,
2444=>134.56529211870634,
2445=>135.22371648265175,
2446=>135.88358818119752,
2447=>136.54490566084314,
2448=>137.20766736468443,
2449=>137.8718717324174,
2450=>138.53751720034165,
2451=>139.20460220136385,
2452=>139.87312516500197,
2453=>140.54308451738837,
2454=>141.21447868127404,
2455=>141.88730607603202,
2456=>142.56156511766096,
2457=>143.2372542187893,
2458=>143.91437178867864,
2459=>144.59291623322758,
2460=>145.27288595497578,
2461=>145.95427935310715,
2462=>146.63709482345405,
2463=>147.32133075850084,
2464=>148.00698554738779,
2465=>148.69405757591483,
2466=>149.38254522654552,
2467=>150.07244687841057,
2468=>150.76376090731173,
2469=>151.45648568572574,
2470=>152.15061958280808,
2471=>152.84616096439663,
2472=>153.543108193016,
2473=>154.2414596278811,
2474=>154.9412136249008,
2475=>155.64236853668194,
2476=>156.3449227125335,
2477=>157.04887449847024,
2478=>157.75422223721625,
2479=>158.4609642682093,
2480=>159.1690989276052,
2481=>159.87862454828064,
2482=>160.58953945983785,
2483=>161.30184198860798,
2484=>162.01553045765593,
2485=>162.73060318678324,
2486=>163.44705849253285,
2487=>164.16489468819293,
2488=>164.88411008380046,
2489=>165.6047029861453,
2490=>166.3266716987746,
2491=>167.05001452199645,
2492=>167.77472975288367,
2493=>168.50081568527878,
2494=>169.2282706097966,
2495=>169.95709281382926,
2496=>170.68728058155034,
2497=>171.41883219391775,
2498=>172.15174592867925,
2499=>172.8860200603757,
2500=>173.62165286034497,
2501=>174.35864259672655,
2502=>175.09698753446548,
2503=>175.8366859353158,
2504=>176.57773605784587,
2505=>177.32013615744142,
2506=>178.0638844863098,
2507=>178.80897929348464,
2508=>179.5554188248293,
2509=>180.30320132304166,
2510=>181.0523250276574,
2511=>181.80278817505564,
2512=>182.5545889984612,
2513=>183.30772572795001,
2514=>184.06219659045303,
2515=>184.8179998097603,
2516=>185.57513360652467,
2517=>186.33359619826751,
2518=>187.09338579938117,
2519=>187.85450062113387,
2520=>188.61693887167428,
2521=>189.38069875603492,
2522=>190.14577847613748,
2523=>190.9121762307957,
2524=>191.67989021572112,
2525=>192.44891862352608,
2526=>193.2192596437285,
2527=>193.99091146275612,
2528=>194.7638722639507,
2529=>195.53814022757228,
2530=>196.31371353080362,
2531=>197.09059034775476,
2532=>197.86876884946616,
2533=>198.64824720391448,
2534=>199.42902357601577,
2535=>200.2110961276303,
2536=>200.9944630175669,
2537=>201.77912240158753,
2538=>202.56507243241072,
2539=>203.35231125971688,
2540=>204.14083703015206,
2541=>204.9306478873326,
2542=>205.7217419718496,
2543=>206.51411742127266,
2544=>207.3077723701556,
2545=>208.10270495003897,
2546=>208.89891328945612,
2547=>209.69639551393686,
2548=>210.49514974601163,
2549=>211.2951741052167,
2550=>212.09646670809752,
2551=>212.89902566821468,
2552=>213.7028490961469,
2553=>214.50793509949597,
2554=>215.31428178289127,
2555=>216.12188724799466,
2556=>216.93074959350395,
2557=>217.740866915158,
2558=>218.55223730574187,
2559=>219.36485885509,
2560=>220.1787296500912,
2561=>220.99384777469334,
2562=>221.81021130990803,
2563=>222.62781833381428,
2564=>223.44666692156466,
2565=>224.26675514538783,
2566=>225.08808107459436,
2567=>225.9106427755811,
2568=>226.73443831183533,
2569=>227.55946574393977,
2570=>228.38572312957672,
2571=>229.21320852353347,
2572=>230.04191997770545,
2573=>230.87185554110226,
2574=>231.70301325985145,
2575=>232.5353911772031,
2576=>233.36898733353496,
2577=>234.20379976635638,
2578=>235.03982651031401,
2579=>235.87706559719493,
2580=>236.71551505593243,
2581=>237.55517291261026,
2582=>238.39603719046727,
2583=>239.2381059099019,
2584=>240.08137708847755,
2585=>240.92584874092648,
2586=>241.77151887915443,
2587=>242.618385512246,
2588=>243.46644664646874,
2589=>244.31570028527818,
2590=>245.16614442932206,
2591=>246.01777707644618,
2592=>246.8705962216976,
2593=>247.7245998573302,
2594=>248.5797859728093,
2595=>249.4361525548166,
2596=>250.29369758725431,
2597=>251.15241905125038,
2598=>252.0123149251636,
2599=>252.8733831845874,
2600=>253.73562180235518,
2601=>254.59902874854532,
2602=>255.46360199048536,
2603=>256.32933949275696,
2604=>257.19623921720165,
2605=>258.06429912292384,
2606=>258.9335171662971,
2607=>259.8038913009681,
2608=>260.67541947786236,
2609=>261.5480996451881,
2610=>262.4219297484415,
2611=>263.2969077304114,
2612=>264.1730315311846,
2613=>265.05029908815004,
2614=>265.92870833600404,
2615=>266.8082572067553,
2616=>267.68894362972924,
2617=>268.57076553157356,
2618=>269.4537208362625,
2619=>270.33780746510206,
2620=>271.22302333673434,
2621=>272.10936636714445,
2622=>272.99683446966236,
2623=>273.8854255549699,
2624=>274.775137531105,
2625=>275.6659683034672,
2626=>276.55791577482097,
2627=>277.4509778453029,
2628=>278.3451524124252,
2629=>279.2404373710811,
2630=>280.13683061354936,
2631=>281.0343300294994,
2632=>281.9329335059979,
2633=>282.83263892751063,
2634=>283.7334441759097,
2635=>284.6353471304781,
2636=>285.5383456679142,
2637=>286.4424376623375,
2638=>287.347620985293,
2639=>288.2538935057564,
2640=>289.1612530901393,
2641=>290.0696976022942,
2642=>290.979224903519,
2643=>291.88983285256285,
2644=>292.80151930563005,
2645=>293.7142821163875,
2646=>294.6281191359665,
2647=>295.54302821296983,
2648=>296.45900719347657,
2649=>297.37605392104683,
2650=>298.2941662367271,
2651=>299.213341979055,
2652=>300.1335789840648,
2653=>301.0548750852923,
2654=>301.9772281137797,
2655=>302.90063589808113,
2656=>303.82509626426764,
2657=>304.7506070359319,
2658=>305.67716603419365,
2659=>306.6047710777059,
2660=>307.5334199826576,
2661=>308.4631105627811,
2662=>309.39384062935585,
2663=>310.32560799121444,
2664=>311.25841045474715,
2665=>312.1922458239076,
2666=>313.1271119002177,
2667=>314.0630064827726,
2668=>314.99992736824635,
2669=>315.9378723508966,
2670=>316.87683922257025,
2671=>317.81682577270766,
2672=>318.7578297883505,
2673=>319.69984905414304,
2674=>320.64288135234045,
2675=>321.58692446281265,
2676=>322.5319761630499,
2677=>323.478034228168,
2678=>324.4250964309136,
2679=>325.37316054166934,
2680=>326.3222243284589,
2681=>327.2722855569529,
2682=>328.2233419904734,
2683=>329.1753913899996,
2684=>330.1284315141725,
2685=>331.0824601193023,
2686=>332.0374749593704,
2687=>332.993473786037,
2688=>333.9504543486456,
2689=>334.9084143942287,
2690=>335.86735166751254,
2691=>336.827263910923,
2692=>337.7881488645905,
2693=>338.7500042663554,
2694=>339.7128278517737,
2695=>340.67661735412156,
2696=>341.64137050440166,
2697=>342.6070850313476,
2698=>343.57375866142934,
2699=>344.5413891188605,
2700=>345.50997412560025,
2701=>346.47951140136144,
2702=>347.4499986636147,
2703=>348.4214336275942,
2704=>349.3938140063033,
2705=>350.3671375105192,
2706=>351.341401848799,
2707=>352.31660472748484,
2708=>353.2927438507092,
2709=>354.26981692040044,
2710=>355.24782163628834,
2711=>356.2267556959085,
2712=>357.20661679461045,
2713=>358.1874026255597,
2714=>359.16911087974506,
2715=>360.1517392459839,
2716=>361.13528541092717,
2717=>362.1197470590653,
2718=>363.1051218727335,
2719=>364.091407532117,
2720=>365.0786017152567,
2721=>366.06670209805486,
2722=>367.05570635427983,
2723=>368.04561215557237,
2724=>369.0364171714509,
2725=>370.02811906931595,
2726=>371.0207155144585,
2727=>372.0142041700618,
2728=>373.0085826972091,
2729=>374.00384875488874,
2730=>374.99999999999966,
2731=>375.99703408735684,
2732=>376.9949486696966,
2733=>377.99374139768264,
2734=>378.99340991991124,
2735=>379.9939518829167,
2736=>380.9953649311771,
2737=>381.9976467071198,
2738=>383.0007948511265,
2739=>384.0048070015407,
2740=>385.0096807946703,
2741=>386.0154138647952,
2742=>387.02200384417245,
2743=>388.02944836304147,
2744=>389.03774504963013,
2745=>390.04689153015994,
2746=>391.05688542885196,
2747=>392.06772436793193,
2748=>393.0794059676365,
2749=>394.0919278462182,
2750=>395.1052876199515,
2751=>396.1194829031383,
2752=>397.1345113081133,
2753=>398.15037044524996,
2754=>399.1670579229661,
2755=>400.18457134772916,
2756=>401.20290832406226,
2757=>402.2220664545498,
2758=>403.2420433398426,
2759=>404.2628365786644,
2760=>405.28444376781664,
2761=>406.30686250218486,
2762=>407.33009037474307,
2763=>408.3541249765625,
2764=>409.3789638968131,
2765=>410.40460472277204,
2766=>411.4310450398284,
2767=>412.4582824314893,
2768=>413.4863144793851,
2769=>414.5151387632756,
2770=>415.5447528610553,
2771=>416.5751543487594,
2772=>417.6063408005692,
2773=>418.6383097888183,
2774=>419.67105888399766,
2775=>420.704585654762,
2776=>421.7388876679344,
2777=>422.77396248851477,
2778=>423.8098076796816,
2779=>424.84642080280076,
2780=>425.8837994174297,
2781=>426.9219410813242,
2782=>427.9608433504432,
2783=>429.00050377895536,
2784=>430.04091991924423,
2785=>431.0820893219142,
2786=>432.1240095357966,
2787=>433.1666781079547,
2788=>434.2100925836903,
2789=>435.2542505065485,
2790=>436.29914941832584,
2791=>437.3447868590727,
2792=>438.39116036710124,
2793=>439.4382674789909,
2794=>440.4861057295939,
2795=>441.5346726520413,
2796=>442.58396577774863,
2797=>443.63398263642165,
2798=>444.6847207560625,
2799=>445.73617766297514,
2800=>446.7883508817714,
2801=>447.8412379353766,
2802=>448.8948363450351,
2803=>449.94914363031825,
2804=>451.00415730912675,
2805=>452.0598748976988,
2806=>453.1162939106157,
2807=>454.17341186080705,
2808=>455.23122625955716,
2809=>456.2897346165108,
2810=>457.3489344396789,
2811=>458.4088232354445,
2812=>459.46939850856864,
2813=>460.53065776219626,
2814=>461.592598497862,
2815=>462.65521821549623,
2816=>463.71851441342994,
2817=>464.7824845884038,
2818=>465.8471262355694,
2819=>466.91243684849866,
2820=>467.9784139191882,
2821=>469.0450549380658,
2822=>470.11235739399615,
2823=>471.18031877428666,
2824=>472.24893656469357,
2825=>473.31820824942776,
2826=>474.38813131116063,
2827=>475.45870323103014,
2828=>476.52992148864655,
2829=>477.60178356209803,
2830=>478.6742869279588,
2831=>479.74742906129154,
2832=>480.8212074356556,
2833=>481.8956195231126,
2834=>482.97066279423217,
2835=>484.0463347180981,
2836=>485.1226327623139,
2837=>486.19955439300935,
2838=>487.277097074846,
2839=>488.3552582710232,
2840=>489.4340354432845,
2841=>490.51342605192286,
2842=>491.59342755578734,
2843=>492.67403741228816,
2844=>493.7552530774051,
2845=>494.83707200568983,
2846=>495.9194916502746,
2847=>497.0025094628772,
2848=>498.0861228938073,
2849=>499.17032939197236,
2850=>500.25512640488364,
2851=>501.3405113786621,
2852=>502.42648175804436,
2853=>503.51303498638913,
2854=>504.60016850568286,
2855=>505.6878797565457,
2856=>506.7761661782374,
2857=>507.8650252086651,
2858=>508.9544542843861,
2859=>510.0444508406165,
2860=>511.13501231123627,
2861=>512.2261361287954,
2862=>513.3178197245201,
2863=>514.4100605283185,
2864=>515.5028559687871,
2865=>516.5962034732166,
2866=>517.6901004675982,
2867=>518.7845443766291,
2868=>519.8795326237193,
2869=>520.9750626309963,
2870=>522.0711318193142,
2871=>523.1677376082562,
2872=>524.2648774161421,
2873=>525.3625486600351,
2874=>526.4607487557471,
2875=>527.559475117845,
2876=>528.6587251596565,
2877=>529.7584962932767,
2878=>530.8587859295737,
2879=>531.9595914781952,
2880=>533.0609103475741,
2881=>534.1627399449349,
2882=>535.2650776762995,
2883=>536.3679209464939,
2884=>537.4712671591537,
2885=>538.5751137167305,
2886=>539.679458020498,
2887=>540.784297470558,
2888=>541.8896294658467,
2889=>542.9954514041408,
2890=>544.1017606820632,
2891=>545.2085546950898,
2892=>546.3158308375552,
2893=>547.4235865026585,
2894=>548.5318190824714,
2895=>549.6405259679415,
2896=>550.7497045488997,
2897=>551.859352214067,
2898=>552.9694663510597,
2899=>554.0800443463963,
2900=>555.1910835855026,
2901=>556.3025814527193,
2902=>557.4145353313068,
2903=>558.5269426034522,
2904=>559.6398006502751,
2905=>560.753106851834,
2906=>561.8668585871321,
2907=>562.9810532341232,
2908=>564.0956881697206,
2909=>565.2107607697985,
2910=>566.3262684092018,
2911=>567.4422084617512,
2912=>568.5585783002491,
2913=>569.6753752964865,
2914=>570.7925968212486,
2915=>571.9102402443208,
2916=>573.0283029344957,
2917=>574.1467822595789,
2918=>575.2656755863947,
2919=>576.384980280793,
2920=>577.5046937076546,
2921=>578.6248132308999,
2922=>579.7453362134916,
2923=>580.8662600174425,
2924=>581.9875820038226,
2925=>583.109299532764,
2926=>584.2314099634677,
2927=>585.3539106542098,
2928=>586.4767989623475,
2929=>587.6000722443255,
2930=>588.723727855682,
2931=>589.8477631510556,
2932=>590.9721754841904,
2933=>592.0969622079434,
2934=>593.2221206742893,
2935=>594.3476482343295,
2936=>595.4735422382947,
2937=>596.5998000355534,
2938=>597.7264189746177,
2939=>598.8533964031494,
2940=>599.9807296679666,
2941=>601.1084161150493,
2942=>602.2364530895463,
2943=>603.364837935781,
2944=>604.493567997258,
2945=>605.6226406166691,
2946=>606.7520531358995,
2947=>607.8818028960336,
2948=>609.0118872373641,
2949=>610.1423034993936,
2950=>611.2730490208443,
2951=>612.404121139663,
2952=>613.5355171930277,
2953=>614.6672345173538,
2954=>615.7992704483003,
2955=>616.9316223207761,
2956=>618.0642874689466,
2957=>619.1972632262391,
2958=>620.3305469253503,
2959=>621.4641358982512,
2960=>622.5980274761948,
2961=>623.7322189897206,
2962=>624.8667077686641,
2963=>626.0014911421591,
2964=>627.1365664386464,
2965=>628.2719309858794,
2966=>629.4075821109307,
2967=>630.5435171401982,
2968=>631.6797333994114,
2969=>632.8162282136378,
2970=>633.952998907289,
2971=>635.0900428041272,
2972=>636.2273572272712,
2973=>637.3649394992033,
2974=>638.5027869417742,
2975=>639.6408968762124,
2976=>640.7792666231267,
2977=>641.9178935025145,
2978=>643.056774833768,
2979=>644.1959079356807,
2980=>645.3352901264526,
2981=>646.4749187236981,
2982=>647.6147910444511,
2983=>648.7549044051717,
2984=>649.8952561217525,
2985=>651.0358435095252,
2986=>652.1766638832664,
2987=>653.3177145572038,
2988=>654.4589928450246,
2989=>655.6004960598783,
2990=>656.7422215143856,
2991=>657.8841665206439,
2992=>659.0263283902339,
2993=>660.1687044342253,
2994=>661.3112919631842,
2995=>662.4540882871783,
2996=>663.5970907157839,
2997=>664.7402965580923,
2998=>665.8837031227155,
2999=>667.0273077177933,
3000=>668.1711076509993,
3001=>669.3151002295461,
3002=>670.4592827601955,
3003=>671.6036525492593,
3004=>672.7482069026098,
3005=>673.8929431256844,
3006=>675.0378585234924,
3007=>676.1829504006214,
3008=>677.3282160612441,
3009=>678.473652809122,
3010=>679.6192579476159,
3011=>680.7650287796889,
3012=>681.910962607916,
3013=>683.0570567344862,
3014=>684.2033084612123,
3015=>685.3497150895354,
3016=>686.4962739205326,
3017=>687.6429822549222,
3018=>688.7898373930708,
3019=>689.9368366349993,
3020=>691.0839772803893,
3021=>692.2312566285893,
3022=>693.3786719786219,
3023=>694.526220629189,
3024=>695.6738998786786,
3025=>696.8217070251709,
3026=>697.9696393664469,
3027=>699.1176941999908,
3028=>700.265868822999,
3029=>701.4141605323861,
3030=>702.5625666247909,
3031=>703.711084396583,
3032=>704.859711143869,
3033=>706.0084441624991,
3034=>707.157280748073,
3035=>708.306218195947,
3036=>709.4552538012397,
3037=>710.6043848588383,
3038=>711.7536086634054,
3039=>712.9029225093865,
3040=>714.0523236910136,
3041=>715.2018095023134,
3042=>716.3513772371136,
3043=>717.5010241890492,
3044=>718.650747651568,
3045=>719.8005449179386,
3046=>720.9504132812552,
3047=>722.1003500344449,
3048=>723.2503524702736,
3049=>724.4004178813526,
3050=>725.5505435601452,
3051=>726.7007267989727,
3052=>727.8509648900199,
3053=>729.001255125345,
3054=>730.1515947968809,
3055=>731.3019811964451,
3056=>732.4524116157452,
3057=>733.6028833463848,
3058=>734.7533936798706,
3059=>735.9039399076181,
3060=>737.0545193209587,
3061=>738.2051292111452,
3062=>739.3557668693588,
3063=>740.5064295867157,
3064=>741.6571146542727,
3065=>742.8078193630333,
3066=>743.9585410039571,
3067=>745.1092768679615,
3068=>746.2600242459312,
3069=>747.4107804287238,
3070=>748.5615427071762,
3071=>749.7123083721109,
3072=>750.8630747143425,
3073=>752.0138390246839,
3074=>753.1645985939529,
3075=>754.3153507129782,
3076=>755.4660926726065,
3077=>756.616821763708,
3078=>757.7675352771828,
3079=>758.9182305039694,
3080=>760.0689047350477,
3081=>761.2195552614473,
3082=>762.370179374254,
3083=>763.5207743646155,
3084=>764.6713375237482,
3085=>765.8218661429433,
3086=>766.9723575135736,
3087=>768.1228089270992,
3088=>769.2732176750745,
3089=>770.4235810491544,
3090=>771.5738963411006,
3091=>772.7241608427878,
3092=>773.8743718462098,
3093=>775.0245266434883,
3094=>776.1746225268753,
3095=>777.3246567887621,
3096=>778.4746267216854,
3097=>779.6245296183329,
3098=>780.7743627715502,
3099=>781.9241234743474,
3100=>783.0738090199051,
3101=>784.2234167015804,
3102=>785.3729438129142,
3103=>786.5223876476368,
3104=>787.6717454996749,
3105=>788.8210146631565,
3106=>789.9701924324206,
3107=>791.1192761020195,
3108=>792.2682629667275,
3109=>793.417150321547,
3110=>794.5659354617144,
3111=>795.7146156827071,
3112=>796.863188280249,
3113=>798.0116505503178,
3114=>799.1599997891509,
3115=>800.3082332932516,
3116=>801.4563483593959,
3117=>802.6043422846383,
3118=>803.7522123663189,
3119=>804.8999559020684,
3120=>806.0475701898176,
3121=>807.1950525277994,
3122=>808.3424002145582,
3123=>809.4896105489552,
3124=>810.6366808301751,
3125=>811.7836083577324,
3126=>812.9303904314775,
3127=>814.0770243516032,
3128=>815.2235074186514,
3129=>816.3698369335186,
3130=>817.5160101974636,
3131=>818.6620245121122,
3132=>819.8078771794643,
3133=>820.9535655019022,
3134=>822.099086782193,
3135=>823.2444383234979,
3136=>824.3896174293776,
3137=>825.5346214037995,
3138=>826.6794475511412,
3139=>827.8240931762009,
3140=>828.9685555842015,
3141=>830.1128320807966,
3142=>831.2569199720781,
3143=>832.400816564581,
3144=>833.5445191652926,
3145=>834.688025081655,
3146=>835.8313316215739,
3147=>836.9744360934246,
3148=>838.1173358060579,
3149=>839.2600280688067,
3150=>840.4025101914924,
3151=>841.544779484431,
3152=>842.6868332584396,
3153=>843.8286688248428,
3154=>844.9702834954785,
3155=>846.1116745827053,
3156=>847.2528393994069,
3157=>848.393775259002,
3158=>849.5344794754463,
3159=>850.6749493632415,
3160=>851.8151822374408,
3161=>852.9551754136556,
3162=>854.0949262080617,
3163=>855.234431937405,
3164=>856.3736899190092,
3165=>857.5126974707803,
3166=>858.6514519112145,
3167=>859.7899505594038,
3168=>860.9281907350422,
3169=>862.0661697584326,
3170=>863.2038849504914,
3171=>864.3413336327587,
3172=>865.4785131274,
3173=>866.6154207572147,
3174=>867.7520538456428,
3175=>868.8884097167703,
3176=>870.024485695336,
3177=>871.1602791067376,
3178=>872.295787277038,
3179=>873.4310075329716,
3180=>874.5659372019508,
3181=>875.7005736120717,
3182=>876.8349140921214,
3183=>877.9689559715824,
3184=>879.1026965806428,
3185=>880.2361332501974,
3186=>881.3692633118577,
3187=>882.5020840979566,
3188=>883.6345929415554,
3189=>884.7667871764496,
3190=>885.8986641371755,
3191=>887.0302211590165,
3192=>888.1614555780087,
3193=>889.2923647309482,
3194=>890.4229459553967,
3195=>891.5531965896877,
3196=>892.6831139729327,
3197=>893.8126954450294,
3198=>894.9419383466645,
3199=>896.0708400193228,
3200=>897.1993978052915,
3201=>898.3276090476681,
3202=>899.4554710903662,
3203=>900.5829812781208,
3204=>901.7101369564955,
3205=>902.8369354718886,
3206=>903.9633741715394,
3207=>905.0894504035339,
3208=>906.2151615168118,
3209=>907.340504861172,
3210=>908.465477787279,
3211=>909.5900776466711,
3212=>910.714301791763,
3213=>911.8381475758542,
3214=>912.9616123531356,
3215=>914.0846934786946,
3216=>915.207388308522,
3217=>916.3296941995179,
3218=>917.4516085094983,
3219=>918.5731285972009,
3220=>919.6942518222916,
3221=>920.8149755453703,
3222=>921.9352971279778,
3223=>923.055213932601,
3224=>924.1747233226814,
3225=>925.2938226626179,
3226=>926.4125093177754,
3227=>927.5307806544902,
3228=>928.6486340400766,
3229=>929.7660668428327,
3230=>930.8830764320469,
3231=>931.9996601780038,
3232=>933.1158154519904,
3233=>934.231539626303,
3234=>935.3468300742521,
3235=>936.4616841701699,
3236=>937.5760992894154,
3237=>938.6900728083808,
3238=>939.8036021044995,
3239=>940.9166845562493,
3240=>942.0293175431599,
3241=>943.1414984458198,
3242=>944.2532246458816,
3243=>945.3644935260681,
3244=>946.4753024701794,
3245=>947.5856488630976,
3246=>948.6955300907944,
3247=>949.8049435403361,
3248=>950.9138865998909,
3249=>952.0223566587339,
3250=>953.1303511072532,
3251=>954.2378673369586,
3252=>955.3449027404839,
3253=>956.4514547115955,
3254=>957.5575206451975,
3255=>958.663097937339,
3256=>959.768183985219,
3257=>960.872776187193,
3258=>961.9768719427793,
3259=>963.080468652665,
3260=>964.1835637187119,
3261=>965.2861545439627,
3262=>966.3882385326475,
3263=>967.4898130901888,
3264=>968.5908756232113,
3265=>969.6914235395407,
3266=>970.7914542482172,
3267=>971.8909651594979,
3268=>972.9899536848638,
3269=>974.0884172370255,
3270=>975.1863532299295,
3271=>976.2837590787644,
3272=>977.3806321999671,
3273=>978.4769700112281,
3274=>979.5727699314982,
3275=>980.6680293809959,
3276=>981.7627457812105,
3277=>982.8569165549102,
3278=>983.9505391261478,
3279=>985.0436109202669,
3280=>986.1361293639077,
3281=>987.2280918850128,
3282=>988.3194959128339,
3283=>989.4103388779374,
3284=>990.5006182122108,
3285=>991.5903313488682,
3286=>992.6794757224568,
3287=>993.7680487688623,
3288=>994.8560479253172,
3289=>995.9434706304031,
3290=>997.0303143240595,
3291=>998.1165764475892,
3292=>999.2022544436637,
3293=>1000.2873457563301,
3294=>1001.3718478310163,
3295=>1002.455758114538,
3296=>1003.5390740551034,
3297=>1004.6217931023205,
3298=>1005.7039127072022,
3299=>1006.7854303221729,
3300=>1007.8663434010741,
3301=>1008.9466493991697,
3302=>1010.0263457731551,
3303=>1011.1054299811585,
3304=>1012.1838994827507,
3305=>1013.261751738949,
3306=>1014.3389842122237,
3307=>1015.415594366505,
3308=>1016.4915796671878,
3309=>1017.5669375811376,
3310=>1018.6416655766977,
3311=>1019.7157611236939,
3312=>1020.7892216934413,
3313=>1021.8620447587491,
3314=>1022.9342277939279,
3315=>1024.0057682747959,
3316=>1025.076663678683,
3317=>1026.1469114844374,
3318=>1027.216509172433,
3319=>1028.2854542245736,
3320=>1029.3537441242995,
3321=>1030.4213763565936,
3322=>1031.488348407987,
3323=>1032.5546577665648,
3324=>1033.620301921973,
3325=>1034.6852783654224,
3326=>1035.749584589697,
3327=>1036.813218089158,
3328=>1037.87617635975,
3329=>1038.9384568990085,
3330=>1040.0000572060637,
3331=>1041.0609747816475,
3332=>1042.1212071280984,
3333=>1043.1807517493687,
3334=>1044.23960615103,
3335=>1045.2977678402785,
3336=>1046.3552343259414,
3337=>1047.4120031184823,
3338=>1048.4680717300075,
3339=>1049.5234376742717,
3340=>1050.578098466684,
3341=>1051.6320516243127,
3342=>1052.685294665894,
3343=>1053.7378251118344,
3344=>1054.7896404842177,
3345=>1055.8407383068125,
3346=>1056.8911161050753,
3347=>1057.940771406159,
3348=>1058.9897017389162,
3349=>1060.0379046339076,
3350=>1061.085377623405,
3351=>1062.1321182413997,
3352=>1063.1781240236069,
3353=>1064.2233925074713,
3354=>1065.267921232174,
3355=>1066.311707738637,
3356=>1067.3547495695311,
3357=>1068.3970442692787,
3358=>1069.4385893840617,
3359=>1070.4793824618264,
3360=>1071.5194210522905,
3361=>1072.5587027069466,
3362=>1073.5972249790705,
3363=>1074.634985423725,
3364=>1075.6719815977672,
3365=>1076.7082110598526,
3366=>1077.7436713704424,
3367=>1078.778360091808,
3368=>1079.8122747880375,
3369=>1080.845413025042,
3370=>1081.8777723705598,
3371=>1082.9093503941626,
3372=>1083.9401446672628,
3373=>1084.9701527631162,
3374=>1085.9993722568308,
3375=>1087.0278007253708,
3376=>1088.0554357475623,
3377=>1089.0822749041,
3378=>1090.1083157775518,
3379=>1091.133555952365,
3380=>1092.157993014872,
3381=>1093.181624553296,
3382=>1094.2044481577566,
3383=>1095.2264614202757,
3384=>1096.2476619347824,
3385=>1097.2680472971197,
3386=>1098.287615105049,
3387=>1099.306362958257,
3388=>1100.3242884583613,
3389=>1101.341389208914,
3390=>1102.35766281541,
3391=>1103.3731068852917,
3392=>1104.3877190279536,
3393=>1105.401496854749,
3394=>1106.4144379789955,
3395=>1107.426540015981,
3396=>1108.4378005829676,
3397=>1109.4482172991998,
3398=>1110.457787785908,
3399=>1111.4665096663148,
3400=>1112.4743805656406,
3401=>1113.4813981111097,
3402=>1114.4875599319548,
3403=>1115.4928636594236,
3404=>1116.497306926784,
3405=>1117.5008873693284,
3406=>1118.5036026243833,
3407=>1119.5054503313095,
3408=>1120.506428131511,
3409=>1121.5065336684397,
3410=>1122.5057645876016,
3411=>1123.5041185365608,
3412=>1124.5015931649468,
3413=>1125.4981861244592,
3414=>1126.4938950688725,
3415=>1127.4887176540433,
3416=>1128.482651537914,
3417=>1129.4756943805205,
3418=>1130.467843843995,
3419=>1131.4590975925735,
3420=>1132.4494532926017,
3421=>1133.4389086125382,
3422=>1134.4274612229617,
3423=>1135.4151087965763,
3424=>1136.4018490082167,
3425=>1137.3876795348535,
3426=>1138.3725980555994,
3427=>1139.3566022517136,
3428=>1140.3396898066085,
3429=>1141.3218584058538,
3430=>1142.3031057371834,
3431=>1143.2834294904994,
3432=>1144.2628273578782,
3433=>1145.2412970335772,
3434=>1146.2188362140378,
3435=>1147.1954425978922,
3436=>1148.1711138859687,
3437=>1149.1458477812969,
3438=>1150.1196419891137,
3439=>1151.0924942168679,
3440=>1152.064402174226,
3441=>1153.0353635730776,
3442=>1154.005376127541,
3443=>1154.9744375539676,
3444=>1155.9425455709488,
3445=>1156.9096978993198,
3446=>1157.8758922621657,
3447=>1158.8411263848286,
3448=>1159.8053979949093,
3449=>1160.768704822275,
3450=>1161.7310445990647,
3451=>1162.6924150596938,
3452=>1163.6528139408597,
3453=>1164.6122389815473,
3454=>1165.5706879230338,
3455=>1166.5281585088949,
3456=>1167.484648485009,
3457=>1168.4401555995637,
3458=>1169.3946776030602,
3459=>1170.3482122483183,
3460=>1171.300757290484,
3461=>1172.252310487031,
3462=>1173.2028695977694,
3463=>1174.1524323848494,
3464=>1175.1009966127663,
3465=>1176.0485600483667,
3466=>1176.995120460853,
3467=>1177.9406756217895,
3468=>1178.8852233051064,
3469=>1179.8287612871063,
3470=>1180.7712873464686,
3471=>1181.7127992642552,
3472=>1182.6532948239148,
3473=>1183.5927718112907,
3474=>1184.5312280146222,
3475=>1185.4686612245528,
3476=>1186.405069234134,
3477=>1187.340449838831,
3478=>1188.274800836528,
3479=>1189.2081200275325,
3480=>1190.1404052145817,
3481=>1191.0716542028472,
3482=>1192.0018647999393,
3483=>1192.9310348159138,
3484=>1193.8591620632758,
3485=>1194.7862443569854,
3486=>1195.7122795144626,
3487=>1196.6372653555936,
3488=>1197.5611997027336,
3489=>1198.4840803807142,
3490=>1199.405905216847,
3491=>1200.3266720409297,
3492=>1201.2463786852504,
3493=>1202.1650229845939,
3494=>1203.0826027762453,
3495=>1203.999115899996,
3496=>1204.9145601981486,
3497=>1205.8289335155223,
3498=>1206.7422336994573,
3499=>1207.6544585998197,
3500=>1208.5656060690085,
3501=>1209.4756739619584,
3502=>1210.3846601361454,
3503=>1211.2925624515924,
3504=>1212.1993787708743,
3505=>1213.1051069591222,
3506=>1214.0097448840293,
3507=>1214.913290415855,
3508=>1215.8157414274312,
3509=>1216.7170957941662,
3510=>1217.61735139405,
3511=>1218.5165061076596,
3512=>1219.4145578181635,
3513=>1220.3115044113265,
3514=>1221.207343775517,
3515=>1222.1020738017078,
3516=>1222.9956923834848,
3517=>1223.88819741705,
3518=>1224.7795868012263,
3519=>1225.6698584374647,
3520=>1226.5590102298465,
3521=>1227.4470400850894,
3522=>1228.3339459125527,
3523=>1229.2197256242418,
3524=>1230.1043771348138,
3525=>1230.9878983615815,
3526=>1231.870287224518,
3527=>1232.7515416462636,
3528=>1233.631659552128,
3529=>1234.5106388700974,
3530=>1235.3884775308381,
3531=>1236.2651734677022,
3532=>1237.1407246167316,
3533=>1238.0151289166636,
3534=>1238.8883843089357,
3535=>1239.760488737689,
3536=>1240.6314401497762,
3537=>1241.5012364947622,
3538=>1242.3698757249338,
3539=>1243.2373557953,
3540=>1244.1036746635991,
3541=>1244.9688302903037,
3542=>1245.8328206386245,
3543=>1246.6956436745158,
3544=>1247.55729736668,
3545=>1248.4177796865717,
3546=>1249.2770886084047,
3547=>1250.1352221091538,
3548=>1250.992178168562,
3549=>1251.8479547691438,
3550=>1252.7025498961902,
3551=>1253.555961537775,
3552=>1254.4081876847563,
3553=>1255.2592263307847,
3554=>1256.109075472306,
3555=>1256.9577331085657,
3556=>1257.8051972416151,
3557=>1258.6514658763156,
3558=>1259.4965370203422,
3559=>1260.3404086841897,
3560=>1261.1830788811767,
3561=>1262.0245456274502,
3562=>1262.86480694199,
3563=>1263.703860846615,
3564=>1264.5417053659858,
3565=>1265.3783385276101,
3566=>1266.2137583618478,
3567=>1267.0479629019148,
3568=>1267.8809501838887,
3569=>1268.7127182467125,
3570=>1269.5432651321994,
3571=>1270.372588885038,
3572=>1271.200687552796,
3573=>1272.0275591859254,
3574=>1272.8532018377668,
3575=>1273.6776135645546,
3576=>1274.500792425421,
3577=>1275.3227364823993,
3578=>1276.1434438004326,
3579=>1276.9629124473734,
3580=>1277.7811404939907,
3581=>1278.5981260139743,
3582=>1279.4138670839397,
3583=>1280.2283617834314,
3584=>1281.0416081949288,
3585=>1281.8536044038497,
3586=>1282.6643484985552,
3587=>1283.4738385703545,
3588=>1284.2820727135086,
3589=>1285.0890490252355,
3590=>1285.8947656057144,
3591=>1286.6992205580905,
3592=>1287.5024119884788,
3593=>1288.3043380059694,
3594=>1289.104996722631,
3595=>1289.904386253516,
3596=>1290.7025047166646,
3597=>1291.49935023311,
3598=>1292.2949209268813,
3599=>1293.08921492501,
3600=>1293.8822303575323,
3601=>1294.673965357495,
3602=>1295.4644180609587,
3603=>1296.2535866070036,
3604=>1297.0414691377327,
3605=>1297.828063798277,
3606=>1298.613368736799,
3607=>1299.3973821044979,
3608=>1300.1801020556131,
3609=>1300.9615267474292,
3610=>1301.7416543402805,
3611=>1302.5204829975546,
3612=>1303.2980108856975,
3613=>1304.0742361742168,
3614=>1304.849157035688,
3615=>1305.622771645756,
3616=>1306.395078183142,
3617=>1307.166074829646,
3618=>1307.9357597701533,
3619=>1308.7041311926355,
3620=>1309.4711872881571,
3621=>1310.23692625088,
3622=>1311.0013462780657,
3623=>1311.7644455700818,
3624=>1312.5262223304046,
3625=>1313.2866747656244,
3626=>1314.0458010854488,
3627=>1314.803599502708,
3628=>1315.5600682333582,
3629=>1316.3152054964858,
3630=>1317.0690095143118,
3631=>1317.8214785121957,
3632=>1318.5726107186413,
3633=>1319.3224043652983,
3634=>1320.0708576869679,
3635=>1320.817968921607,
3636=>1321.5637363103315,
3637=>1322.3081580974222,
3638=>1323.0512325303266,
3639=>1323.792957859665,
3640=>1324.5333323392333,
3641=>1325.272354226008,
3642=>1326.0100217801496,
3643=>1326.7463332650075,
3644=>1327.4812869471225,
3645=>1328.2148810962344,
3646=>1328.9471139852808,
3647=>1329.6779838904058,
3648=>1330.407489090962,
3649=>1331.135627869515,
3650=>1331.862398511846,
3651=>1332.587799306959,
3652=>1333.3118285470814,
3653=>1334.0344845276709,
3654=>1334.755765547417,
3655=>1335.4756699082468,
3656=>1336.1941959153291,
3657=>1336.9113418770762,
3658=>1337.6271061051505,
3659=>1338.3414869144667,
3660=>1339.0544826231967,
3661=>1339.766091552773,
3662=>1340.4763120278935,
3663=>1341.1851423765247,
3664=>1341.8925809299049,
3665=>1342.59862602255,
3666=>1343.3032759922562,
3667=>1344.006529180104,
3668=>1344.7083839304623,
3669=>1345.4088385909934,
3670=>1346.1078915126536,
3671=>1346.8055410497009,
3672=>1347.5017855596961,
3673=>1348.196623403509,
3674=>1348.8900529453203,
3675=>1349.582072552626,
3676=>1350.2726805962416,
3677=>1350.9618754503063,
3678=>1351.6496554922858,
3679=>1352.3360191029765,
3680=>1353.0209646665098,
3681=>1353.7044905703547,
3682=>1354.3865952053243,
3683=>1355.0672769655753,
3684=>1355.7465342486164,
3685=>1356.4243654553084,
3686=>1357.1007689898697,
3687=>1357.7757432598805,
3688=>1358.4492866762848,
3689=>1359.121397653396,
3690=>1359.7920746088994,
3691=>1360.4613159638566,
3692=>1361.1291201427089,
3693=>1361.7954855732805,
3694=>1362.460410686784,
3695=>1363.123893917821,
3696=>1363.7859337043901,
3697=>1364.446528487886,
3698=>1365.1056767131063,
3699=>1365.763376828254,
3700=>1366.4196272849413,
3701=>1367.0744265381927,
3702=>1367.7277730464502,
3703=>1368.379665271575,
3704=>1369.0301016788528,
3705=>1369.6790807369962,
3706=>1370.3266009181489,
3707=>1370.9726606978888,
3708=>1371.6172585552322,
3709=>1372.2603929726379,
3710=>1372.9020624360087,
3711=>1373.542265434697,
3712=>1374.1810004615072,
3713=>1374.8182660127004,
3714=>1375.4540605879965,
3715=>1376.0883826905788,
3716=>1376.7212308270964,
3717=>1377.3526035076702,
3718=>1377.9824992458925,
3719=>1378.6109165588346,
3720=>1379.2378539670472,
3721=>1379.8633099945653,
3722=>1380.4872831689113,
3723=>1381.1097720210998,
3724=>1381.7307750856385,
3725=>1382.350290900533,
3726=>1382.9683180072914,
3727=>1383.584854950925,
3728=>1384.199900279955,
3729=>1384.813452546413,
3730=>1385.4255103058458,
3731=>1386.0360721173195,
3732=>1386.645136543421,
3733=>1387.2527021502624,
3734=>1387.8587675074857,
3735=>1388.463331188263,
3736=>1389.0663917693037,
3737=>1389.6679478308542,
3738=>1390.2679979567038,
3739=>1390.8665407341869,
3740=>1391.4635747541865,
3741=>1392.0590986111374,
3742=>1392.6531109030304,
3743=>1393.245610231414,
3744=>1393.8365952013996,
3745=>1394.4260644216624,
3746=>1395.0140165044477,
3747=>1395.600450065571,
3748=>1396.1853637244235,
3749=>1396.7687561039752,
3750=>1397.3506258307764,
3751=>1397.9309715349627,
3752=>1398.509791850258,
3753=>1399.087085413976,
3754=>1399.662850867026,
3755=>1400.2370868539151,
3756=>1400.8097920227497,
3757=>1401.3809650252415,
3758=>1401.9506045167086,
3759=>1402.5187091560792,
3760=>1403.085277605896,
3761=>1403.6503085323166,
3762=>1404.213800605119,
3763=>1404.7757524977058,
3764=>1405.3361628871025,
3765=>1405.8950304539662,
3766=>1406.4523538825847,
3767=>1407.0081318608813,
3768=>1407.5623630804184,
3769=>1408.115046236399,
3770=>1408.666180027671,
3771=>1409.2157631567306,
3772=>1409.7637943297232,
3773=>1410.3102722564486,
3774=>1410.8551956503634,
3775=>1411.398563228584,
3776=>1411.9403737118898,
3777=>1412.4806258247252,
3778=>1413.019318295204,
3779=>1413.5564498551112,
3780=>1414.0920192399076,
3781=>1414.6260251887306,
3782=>1415.1584664443992,
3783=>1415.6893417534156,
3784=>1416.218649865969,
3785=>1416.7463895359372,
3786=>1417.2725595208913,
3787=>1417.7971585820987,
3788=>1418.3201854845233,
3789=>1418.8416389968313,
3790=>1419.3615178913929,
3791=>1419.8798209442853,
3792=>1420.3965469352956,
3793=>1420.9116946479237,
3794=>1421.425262869385,
3795=>1421.9372503906138,
3796=>1422.4476560062658,
3797=>1422.95647851472,
3798=>1423.4637167180833,
3799=>1423.969369422192,
3800=>1424.4734354366158,
3801=>1424.975913574659,
3802=>1425.4768026533643,
3803=>1425.9761014935161,
3804=>1426.4738089196417,
3805=>1426.969923760015,
3806=>1427.4644448466604,
3807=>1427.9573710153531,
3808=>1428.4487011056242,
3809=>1428.9384339607611,
3810=>1429.4265684278125,
3811=>1429.91310335759,
3812=>1430.3980376046707,
3813=>1430.881370027399,
3814=>1431.3630994878931,
3815=>1431.8432248520426,
3816=>1432.3217449895142,
3817=>1432.7986587737541,
3818=>1433.2739650819894,
3819=>1433.7476627952328,
3820=>1434.2197507982828,
3821=>1434.6902279797287,
3822=>1435.1590932319507,
3823=>1435.6263454511252,
3824=>1436.0919835372256,
3825=>1436.5560063940247,
3826=>1437.0184129290992,
3827=>1437.47920205383,
3828=>1437.9383726834067,
3829=>1438.3959237368279,
3830=>1438.8518541369062,
3831=>1439.3061628102696,
3832=>1439.7588486873635,
3833=>1440.2099107024537,
3834=>1440.6593477936296,
3835=>1441.1071589028056,
3836=>1441.5533429757243,
3837=>1441.9978989619585,
3838=>1442.4408258149142,
3839=>1442.8821224918327,
3840=>1443.3217879537924,
3841=>1443.7598211657134,
3842=>1444.1962210963577,
3843=>1444.6309867183322,
3844=>1445.0641170080921,
3845=>1445.4956109459415,
3846=>1445.9254675160382,
3847=>1446.3536857063937,
3848=>1446.7802645088768,
3849=>1447.2052029192168,
3850=>1447.6284999370037,
3851=>1448.050154565692,
3852=>1448.4701658126037,
3853=>1448.888532688928,
3854=>1449.305254209727,
3855=>1449.720329393936,
3856=>1450.1337572643654,
3857=>1450.5455368477042,
3858=>1450.9556671745224,
3859=>1451.3641472792722,
3860=>1451.7709762002908,
3861=>1452.1761529798027,
3862=>1452.5796766639228,
3863=>1452.9815463026562,
3864=>1453.3817609499033,
3865=>1453.7803196634604,
3866=>1454.1772215050223,
3867=>1454.5724655401843,
3868=>1454.966050838445,
3869=>1455.3579764732071,
3870=>1455.7482415217821,
3871=>1456.1368450653897,
3872=>1456.5237861891615,
3873=>1456.909063982143,
3874=>1457.2926775372953,
3875=>1457.674625951498,
3876=>1458.0549083255505,
3877=>1458.4335237641744,
3878=>1458.8104713760158,
3879=>1459.1857502736477,
3880=>1459.5593595735709,
3881=>1459.9312983962172,
3882=>1460.3015658659513,
3883=>1460.6701611110725,
3884=>1461.0370832638166,
3885=>1461.4023314603592,
3886=>1461.7659048408154,
3887=>1462.1278025492447,
3888=>1462.4880237336506,
3889=>1462.8465675459838,
3890=>1463.203433142144,
3891=>1463.5586196819818,
3892=>1463.912126329301,
3893=>1464.2639522518589,
3894=>1464.614096621372,
3895=>1464.9625586135141,
3896=>1465.3093374079197,
3897=>1465.654432188186,
3898=>1465.9978421418755,
3899=>1466.3395664605164,
3900=>1466.6796043396055,
3901=>1467.01795497861,
3902=>1467.3546175809697,
3903=>1467.6895913540975,
3904=>1468.0228755093826,
3905=>1468.354469262193,
3906=>1468.6843718318746,
3907=>1469.012582441756,
3908=>1469.3391003191484,
3909=>1469.6639246953487,
3910=>1469.9870548056401,
3911=>1470.3084898892953,
3912=>1470.6282291895766,
3913=>1470.9462719537391,
3914=>1471.2626174330321,
3915=>1471.5772648827005,
3916=>1471.8902135619865,
3917=>1472.2014627341323,
3918=>1472.5110116663805,
3919=>1472.818859629977,
3920=>1473.1250059001718,
3921=>1473.4294497562214,
3922=>1473.7321904813898,
3923=>1474.0332273629513,
3924=>1474.332559692191,
3925=>1474.630186764406,
3926=>1474.9261078789104,
3927=>1475.2203223390322,
3928=>1475.5128294521185,
3929=>1475.8036285295354,
3930=>1476.0927188866706,
3931=>1476.3800998429338,
3932=>1476.66577072176,
3933=>1476.9497308506097,
3934=>1477.2319795609706,
3935=>1477.5125161883602,
3936=>1477.791340072326,
3937=>1478.0684505564477,
3938=>1478.3438469883397,
3939=>1478.6175287196506,
3940=>1478.8894951060665,
3941=>1479.1597455073115,
3942=>1479.4282792871495,
3943=>1479.6950958133864,
3944=>1479.9601944578699,
3945=>1480.223574596493,
3946=>1480.4852356091942,
3947=>1480.7451768799588,
3948=>1481.003397796821,
3949=>1481.2598977518653,
3950=>1481.514676141228,
3951=>1481.7677323650978,
3952=>1482.0190658277184,
3953=>1482.2686759373887,
3954=>1482.5165621064652,
3955=>1482.762723751363,
3956=>1483.0071602925568,
3957=>1483.2498711545827,
3958=>1483.4908557660403,
3959=>1483.7301135595922,
3960=>1483.9676439719665,
3961=>1484.2034464439582,
3962=>1484.4375204204307,
3963=>1484.6698653503158,
3964=>1484.9004806866164,
3965=>1485.1293658864079,
3966=>1485.3565204108374,
3967=>1485.581943725128,
3968=>1485.805635298577,
3969=>1486.02759460456,
3970=>1486.2478211205303,
3971=>1486.4663143280197,
3972=>1486.683073712642,
3973=>1486.8980987640925,
3974=>1487.111388976149,
3975=>1487.3229438466742,
3976=>1487.5327628776154,
3977=>1487.7408455750074,
3978=>1487.9471914489723,
3979=>1488.1518000137207,
3980=>1488.3546707875544,
3981=>1488.555803292865,
3982=>1488.7551970561376,
3983=>1488.9528516079502,
3984=>1489.1487664829751,
3985=>1489.3429412199807,
3986=>1489.5353753618317,
3987=>1489.726068455491,
3988=>1489.9150200520203,
3989=>1490.1022297065806,
3990=>1490.2876969784347,
3991=>1490.4714214309467,
3992=>1490.6534026315844,
3993=>1490.833640151919,
3994=>1491.0121335676272,
3995=>1491.1888824584917,
3996=>1491.3638864084019,
3997=>1491.5371450053553,
3998=>1491.7086578414592,
3999=>1491.8784245129295,
4000=>1492.046444620094,
4001=>1492.212717767392,
4002=>1492.3772435633757,
4003=>1492.5400216207108,
4004=>1492.7010515561778,
4005=>1492.8603329906723,
4006=>1493.017865549207,
4007=>1493.1736488609115,
4008=>1493.3276825590333,
4009=>1493.4799662809394,
4010=>1493.6304996681163,
4011=>1493.7792823661714,
4012=>1493.9263140248338,
4013=>1494.0715942979546,
4014=>1494.2151228435087,
4015=>1494.356899323594,
4016=>1494.4969234044343,
4017=>1494.635194756378,
4018=>1494.7717130539006,
4019=>1494.9064779756045,
4020=>1495.03948920422,
4021=>1495.1707464266055,
4022=>1495.3002493337497,
4023=>1495.4279976207708,
4024=>1495.5539909869176,
4025=>1495.6782291355707,
4026=>1495.8007117742436,
4027=>1495.9214386145816,
4028=>1496.040409372364,
4029=>1496.1576237675042,
4030=>1496.2730815240511,
4031=>1496.3867823701885,
4032=>1496.4987260382363,
4033=>1496.6089122646524,
4034=>1496.7173407900307,
4035=>1496.8240113591037,
4036=>1496.9289237207431,
4037=>1497.032077627959,
4038=>1497.1334728379022,
4039=>1497.233109111863,
4040=>1497.3309862152732,
4041=>1497.427103917706,
4042=>1497.5214619928765,
4043=>1497.6140602186433,
4044=>1497.7048983770064,
4045=>1497.7939762541114,
4046=>1497.8812936402464,
4047=>1497.9668503298449,
4048=>1498.0506461214854,
4049=>1498.1326808178924,
4050=>1498.2129542259356,
4051=>1498.291466156632,
4052=>1498.3682164251447,
4053=>1498.4432048507852,
4054=>1498.5164312570118,
4055=>1498.5878954714321,
4056=>1498.6575973258014,
4057=>1498.7255366560244,
4058=>1498.7917133021551,
4059=>1498.856127108398,
4060=>1498.9187779231065,
4061=>1498.9796655987852,
4062=>1499.0387899920897,
4063=>1499.0961509638269,
4064=>1499.1517483789548,
4065=>1499.205582106583,
4066=>1499.257652019974,
4067=>1499.3079579965429,
4068=>1499.3564999178561,
4069=>1499.4032776696345,
4070=>1499.4482911417517,
4071=>1499.491540228235,
4072=>1499.5330248272653,
4073=>1499.5727448411776,
4074=>1499.6107001764613,
4075=>1499.6468907437602,
4076=>1499.6813164578728,
4077=>1499.7139772377525,
4078=>1499.7448730065078,
4079=>1499.7740036914024,
4080=>1499.8013692238555,
4081=>1499.8269695394422,
4082=>1499.8508045778926,
4083=>1499.8728742830936,
4084=>1499.893178603087,
4085=>1499.9117174900723,
4086=>1499.928490900404,
4087=>1499.9434987945933,
4088=>1499.9567411373077,
4089=>1499.9682178973721,
4090=>1499.9779290477668,
4091=>1499.9858745656297,
4092=>1499.992054432255,
4093=>1499.9964686330936,
4094=>1499.999117157754,
4095=>1500.0
    );

signal lut_sig : unsigned(15 downto 0);

begin 
    cos <= STD_LOGIC_VECTOR(lut_sig);
    process (address)
            begin
                case address is
                   when x"000" => lut_sig <= to_unsigned(integer(my_cos(0)),16);
when x"001" => lut_sig <= to_unsigned(integer(my_cos(1)),16);
when x"002" => lut_sig <= to_unsigned(integer(my_cos(2)),16);
when x"003" => lut_sig <= to_unsigned(integer(my_cos(3)),16);
when x"004" => lut_sig <= to_unsigned(integer(my_cos(4)),16);
when x"005" => lut_sig <= to_unsigned(integer(my_cos(5)),16);
when x"006" => lut_sig <= to_unsigned(integer(my_cos(6)),16);
when x"007" => lut_sig <= to_unsigned(integer(my_cos(7)),16);
when x"008" => lut_sig <= to_unsigned(integer(my_cos(8)),16);
when x"009" => lut_sig <= to_unsigned(integer(my_cos(9)),16);
when x"00a" => lut_sig <= to_unsigned(integer(my_cos(10)),16);
when x"00b" => lut_sig <= to_unsigned(integer(my_cos(11)),16);
when x"00c" => lut_sig <= to_unsigned(integer(my_cos(12)),16);
when x"00d" => lut_sig <= to_unsigned(integer(my_cos(13)),16);
when x"00e" => lut_sig <= to_unsigned(integer(my_cos(14)),16);
when x"00f" => lut_sig <= to_unsigned(integer(my_cos(15)),16);
when x"010" => lut_sig <= to_unsigned(integer(my_cos(16)),16);
when x"011" => lut_sig <= to_unsigned(integer(my_cos(17)),16);
when x"012" => lut_sig <= to_unsigned(integer(my_cos(18)),16);
when x"013" => lut_sig <= to_unsigned(integer(my_cos(19)),16);
when x"014" => lut_sig <= to_unsigned(integer(my_cos(20)),16);
when x"015" => lut_sig <= to_unsigned(integer(my_cos(21)),16);
when x"016" => lut_sig <= to_unsigned(integer(my_cos(22)),16);
when x"017" => lut_sig <= to_unsigned(integer(my_cos(23)),16);
when x"018" => lut_sig <= to_unsigned(integer(my_cos(24)),16);
when x"019" => lut_sig <= to_unsigned(integer(my_cos(25)),16);
when x"01a" => lut_sig <= to_unsigned(integer(my_cos(26)),16);
when x"01b" => lut_sig <= to_unsigned(integer(my_cos(27)),16);
when x"01c" => lut_sig <= to_unsigned(integer(my_cos(28)),16);
when x"01d" => lut_sig <= to_unsigned(integer(my_cos(29)),16);
when x"01e" => lut_sig <= to_unsigned(integer(my_cos(30)),16);
when x"01f" => lut_sig <= to_unsigned(integer(my_cos(31)),16);
when x"020" => lut_sig <= to_unsigned(integer(my_cos(32)),16);
when x"021" => lut_sig <= to_unsigned(integer(my_cos(33)),16);
when x"022" => lut_sig <= to_unsigned(integer(my_cos(34)),16);
when x"023" => lut_sig <= to_unsigned(integer(my_cos(35)),16);
when x"024" => lut_sig <= to_unsigned(integer(my_cos(36)),16);
when x"025" => lut_sig <= to_unsigned(integer(my_cos(37)),16);
when x"026" => lut_sig <= to_unsigned(integer(my_cos(38)),16);
when x"027" => lut_sig <= to_unsigned(integer(my_cos(39)),16);
when x"028" => lut_sig <= to_unsigned(integer(my_cos(40)),16);
when x"029" => lut_sig <= to_unsigned(integer(my_cos(41)),16);
when x"02a" => lut_sig <= to_unsigned(integer(my_cos(42)),16);
when x"02b" => lut_sig <= to_unsigned(integer(my_cos(43)),16);
when x"02c" => lut_sig <= to_unsigned(integer(my_cos(44)),16);
when x"02d" => lut_sig <= to_unsigned(integer(my_cos(45)),16);
when x"02e" => lut_sig <= to_unsigned(integer(my_cos(46)),16);
when x"02f" => lut_sig <= to_unsigned(integer(my_cos(47)),16);
when x"030" => lut_sig <= to_unsigned(integer(my_cos(48)),16);
when x"031" => lut_sig <= to_unsigned(integer(my_cos(49)),16);
when x"032" => lut_sig <= to_unsigned(integer(my_cos(50)),16);
when x"033" => lut_sig <= to_unsigned(integer(my_cos(51)),16);
when x"034" => lut_sig <= to_unsigned(integer(my_cos(52)),16);
when x"035" => lut_sig <= to_unsigned(integer(my_cos(53)),16);
when x"036" => lut_sig <= to_unsigned(integer(my_cos(54)),16);
when x"037" => lut_sig <= to_unsigned(integer(my_cos(55)),16);
when x"038" => lut_sig <= to_unsigned(integer(my_cos(56)),16);
when x"039" => lut_sig <= to_unsigned(integer(my_cos(57)),16);
when x"03a" => lut_sig <= to_unsigned(integer(my_cos(58)),16);
when x"03b" => lut_sig <= to_unsigned(integer(my_cos(59)),16);
when x"03c" => lut_sig <= to_unsigned(integer(my_cos(60)),16);
when x"03d" => lut_sig <= to_unsigned(integer(my_cos(61)),16);
when x"03e" => lut_sig <= to_unsigned(integer(my_cos(62)),16);
when x"03f" => lut_sig <= to_unsigned(integer(my_cos(63)),16);
when x"040" => lut_sig <= to_unsigned(integer(my_cos(64)),16);
when x"041" => lut_sig <= to_unsigned(integer(my_cos(65)),16);
when x"042" => lut_sig <= to_unsigned(integer(my_cos(66)),16);
when x"043" => lut_sig <= to_unsigned(integer(my_cos(67)),16);
when x"044" => lut_sig <= to_unsigned(integer(my_cos(68)),16);
when x"045" => lut_sig <= to_unsigned(integer(my_cos(69)),16);
when x"046" => lut_sig <= to_unsigned(integer(my_cos(70)),16);
when x"047" => lut_sig <= to_unsigned(integer(my_cos(71)),16);
when x"048" => lut_sig <= to_unsigned(integer(my_cos(72)),16);
when x"049" => lut_sig <= to_unsigned(integer(my_cos(73)),16);
when x"04a" => lut_sig <= to_unsigned(integer(my_cos(74)),16);
when x"04b" => lut_sig <= to_unsigned(integer(my_cos(75)),16);
when x"04c" => lut_sig <= to_unsigned(integer(my_cos(76)),16);
when x"04d" => lut_sig <= to_unsigned(integer(my_cos(77)),16);
when x"04e" => lut_sig <= to_unsigned(integer(my_cos(78)),16);
when x"04f" => lut_sig <= to_unsigned(integer(my_cos(79)),16);
when x"050" => lut_sig <= to_unsigned(integer(my_cos(80)),16);
when x"051" => lut_sig <= to_unsigned(integer(my_cos(81)),16);
when x"052" => lut_sig <= to_unsigned(integer(my_cos(82)),16);
when x"053" => lut_sig <= to_unsigned(integer(my_cos(83)),16);
when x"054" => lut_sig <= to_unsigned(integer(my_cos(84)),16);
when x"055" => lut_sig <= to_unsigned(integer(my_cos(85)),16);
when x"056" => lut_sig <= to_unsigned(integer(my_cos(86)),16);
when x"057" => lut_sig <= to_unsigned(integer(my_cos(87)),16);
when x"058" => lut_sig <= to_unsigned(integer(my_cos(88)),16);
when x"059" => lut_sig <= to_unsigned(integer(my_cos(89)),16);
when x"05a" => lut_sig <= to_unsigned(integer(my_cos(90)),16);
when x"05b" => lut_sig <= to_unsigned(integer(my_cos(91)),16);
when x"05c" => lut_sig <= to_unsigned(integer(my_cos(92)),16);
when x"05d" => lut_sig <= to_unsigned(integer(my_cos(93)),16);
when x"05e" => lut_sig <= to_unsigned(integer(my_cos(94)),16);
when x"05f" => lut_sig <= to_unsigned(integer(my_cos(95)),16);
when x"060" => lut_sig <= to_unsigned(integer(my_cos(96)),16);
when x"061" => lut_sig <= to_unsigned(integer(my_cos(97)),16);
when x"062" => lut_sig <= to_unsigned(integer(my_cos(98)),16);
when x"063" => lut_sig <= to_unsigned(integer(my_cos(99)),16);
when x"064" => lut_sig <= to_unsigned(integer(my_cos(100)),16);
when x"065" => lut_sig <= to_unsigned(integer(my_cos(101)),16);
when x"066" => lut_sig <= to_unsigned(integer(my_cos(102)),16);
when x"067" => lut_sig <= to_unsigned(integer(my_cos(103)),16);
when x"068" => lut_sig <= to_unsigned(integer(my_cos(104)),16);
when x"069" => lut_sig <= to_unsigned(integer(my_cos(105)),16);
when x"06a" => lut_sig <= to_unsigned(integer(my_cos(106)),16);
when x"06b" => lut_sig <= to_unsigned(integer(my_cos(107)),16);
when x"06c" => lut_sig <= to_unsigned(integer(my_cos(108)),16);
when x"06d" => lut_sig <= to_unsigned(integer(my_cos(109)),16);
when x"06e" => lut_sig <= to_unsigned(integer(my_cos(110)),16);
when x"06f" => lut_sig <= to_unsigned(integer(my_cos(111)),16);
when x"070" => lut_sig <= to_unsigned(integer(my_cos(112)),16);
when x"071" => lut_sig <= to_unsigned(integer(my_cos(113)),16);
when x"072" => lut_sig <= to_unsigned(integer(my_cos(114)),16);
when x"073" => lut_sig <= to_unsigned(integer(my_cos(115)),16);
when x"074" => lut_sig <= to_unsigned(integer(my_cos(116)),16);
when x"075" => lut_sig <= to_unsigned(integer(my_cos(117)),16);
when x"076" => lut_sig <= to_unsigned(integer(my_cos(118)),16);
when x"077" => lut_sig <= to_unsigned(integer(my_cos(119)),16);
when x"078" => lut_sig <= to_unsigned(integer(my_cos(120)),16);
when x"079" => lut_sig <= to_unsigned(integer(my_cos(121)),16);
when x"07a" => lut_sig <= to_unsigned(integer(my_cos(122)),16);
when x"07b" => lut_sig <= to_unsigned(integer(my_cos(123)),16);
when x"07c" => lut_sig <= to_unsigned(integer(my_cos(124)),16);
when x"07d" => lut_sig <= to_unsigned(integer(my_cos(125)),16);
when x"07e" => lut_sig <= to_unsigned(integer(my_cos(126)),16);
when x"07f" => lut_sig <= to_unsigned(integer(my_cos(127)),16);
when x"080" => lut_sig <= to_unsigned(integer(my_cos(128)),16);
when x"081" => lut_sig <= to_unsigned(integer(my_cos(129)),16);
when x"082" => lut_sig <= to_unsigned(integer(my_cos(130)),16);
when x"083" => lut_sig <= to_unsigned(integer(my_cos(131)),16);
when x"084" => lut_sig <= to_unsigned(integer(my_cos(132)),16);
when x"085" => lut_sig <= to_unsigned(integer(my_cos(133)),16);
when x"086" => lut_sig <= to_unsigned(integer(my_cos(134)),16);
when x"087" => lut_sig <= to_unsigned(integer(my_cos(135)),16);
when x"088" => lut_sig <= to_unsigned(integer(my_cos(136)),16);
when x"089" => lut_sig <= to_unsigned(integer(my_cos(137)),16);
when x"08a" => lut_sig <= to_unsigned(integer(my_cos(138)),16);
when x"08b" => lut_sig <= to_unsigned(integer(my_cos(139)),16);
when x"08c" => lut_sig <= to_unsigned(integer(my_cos(140)),16);
when x"08d" => lut_sig <= to_unsigned(integer(my_cos(141)),16);
when x"08e" => lut_sig <= to_unsigned(integer(my_cos(142)),16);
when x"08f" => lut_sig <= to_unsigned(integer(my_cos(143)),16);
when x"090" => lut_sig <= to_unsigned(integer(my_cos(144)),16);
when x"091" => lut_sig <= to_unsigned(integer(my_cos(145)),16);
when x"092" => lut_sig <= to_unsigned(integer(my_cos(146)),16);
when x"093" => lut_sig <= to_unsigned(integer(my_cos(147)),16);
when x"094" => lut_sig <= to_unsigned(integer(my_cos(148)),16);
when x"095" => lut_sig <= to_unsigned(integer(my_cos(149)),16);
when x"096" => lut_sig <= to_unsigned(integer(my_cos(150)),16);
when x"097" => lut_sig <= to_unsigned(integer(my_cos(151)),16);
when x"098" => lut_sig <= to_unsigned(integer(my_cos(152)),16);
when x"099" => lut_sig <= to_unsigned(integer(my_cos(153)),16);
when x"09a" => lut_sig <= to_unsigned(integer(my_cos(154)),16);
when x"09b" => lut_sig <= to_unsigned(integer(my_cos(155)),16);
when x"09c" => lut_sig <= to_unsigned(integer(my_cos(156)),16);
when x"09d" => lut_sig <= to_unsigned(integer(my_cos(157)),16);
when x"09e" => lut_sig <= to_unsigned(integer(my_cos(158)),16);
when x"09f" => lut_sig <= to_unsigned(integer(my_cos(159)),16);
when x"0a0" => lut_sig <= to_unsigned(integer(my_cos(160)),16);
when x"0a1" => lut_sig <= to_unsigned(integer(my_cos(161)),16);
when x"0a2" => lut_sig <= to_unsigned(integer(my_cos(162)),16);
when x"0a3" => lut_sig <= to_unsigned(integer(my_cos(163)),16);
when x"0a4" => lut_sig <= to_unsigned(integer(my_cos(164)),16);
when x"0a5" => lut_sig <= to_unsigned(integer(my_cos(165)),16);
when x"0a6" => lut_sig <= to_unsigned(integer(my_cos(166)),16);
when x"0a7" => lut_sig <= to_unsigned(integer(my_cos(167)),16);
when x"0a8" => lut_sig <= to_unsigned(integer(my_cos(168)),16);
when x"0a9" => lut_sig <= to_unsigned(integer(my_cos(169)),16);
when x"0aa" => lut_sig <= to_unsigned(integer(my_cos(170)),16);
when x"0ab" => lut_sig <= to_unsigned(integer(my_cos(171)),16);
when x"0ac" => lut_sig <= to_unsigned(integer(my_cos(172)),16);
when x"0ad" => lut_sig <= to_unsigned(integer(my_cos(173)),16);
when x"0ae" => lut_sig <= to_unsigned(integer(my_cos(174)),16);
when x"0af" => lut_sig <= to_unsigned(integer(my_cos(175)),16);
when x"0b0" => lut_sig <= to_unsigned(integer(my_cos(176)),16);
when x"0b1" => lut_sig <= to_unsigned(integer(my_cos(177)),16);
when x"0b2" => lut_sig <= to_unsigned(integer(my_cos(178)),16);
when x"0b3" => lut_sig <= to_unsigned(integer(my_cos(179)),16);
when x"0b4" => lut_sig <= to_unsigned(integer(my_cos(180)),16);
when x"0b5" => lut_sig <= to_unsigned(integer(my_cos(181)),16);
when x"0b6" => lut_sig <= to_unsigned(integer(my_cos(182)),16);
when x"0b7" => lut_sig <= to_unsigned(integer(my_cos(183)),16);
when x"0b8" => lut_sig <= to_unsigned(integer(my_cos(184)),16);
when x"0b9" => lut_sig <= to_unsigned(integer(my_cos(185)),16);
when x"0ba" => lut_sig <= to_unsigned(integer(my_cos(186)),16);
when x"0bb" => lut_sig <= to_unsigned(integer(my_cos(187)),16);
when x"0bc" => lut_sig <= to_unsigned(integer(my_cos(188)),16);
when x"0bd" => lut_sig <= to_unsigned(integer(my_cos(189)),16);
when x"0be" => lut_sig <= to_unsigned(integer(my_cos(190)),16);
when x"0bf" => lut_sig <= to_unsigned(integer(my_cos(191)),16);
when x"0c0" => lut_sig <= to_unsigned(integer(my_cos(192)),16);
when x"0c1" => lut_sig <= to_unsigned(integer(my_cos(193)),16);
when x"0c2" => lut_sig <= to_unsigned(integer(my_cos(194)),16);
when x"0c3" => lut_sig <= to_unsigned(integer(my_cos(195)),16);
when x"0c4" => lut_sig <= to_unsigned(integer(my_cos(196)),16);
when x"0c5" => lut_sig <= to_unsigned(integer(my_cos(197)),16);
when x"0c6" => lut_sig <= to_unsigned(integer(my_cos(198)),16);
when x"0c7" => lut_sig <= to_unsigned(integer(my_cos(199)),16);
when x"0c8" => lut_sig <= to_unsigned(integer(my_cos(200)),16);
when x"0c9" => lut_sig <= to_unsigned(integer(my_cos(201)),16);
when x"0ca" => lut_sig <= to_unsigned(integer(my_cos(202)),16);
when x"0cb" => lut_sig <= to_unsigned(integer(my_cos(203)),16);
when x"0cc" => lut_sig <= to_unsigned(integer(my_cos(204)),16);
when x"0cd" => lut_sig <= to_unsigned(integer(my_cos(205)),16);
when x"0ce" => lut_sig <= to_unsigned(integer(my_cos(206)),16);
when x"0cf" => lut_sig <= to_unsigned(integer(my_cos(207)),16);
when x"0d0" => lut_sig <= to_unsigned(integer(my_cos(208)),16);
when x"0d1" => lut_sig <= to_unsigned(integer(my_cos(209)),16);
when x"0d2" => lut_sig <= to_unsigned(integer(my_cos(210)),16);
when x"0d3" => lut_sig <= to_unsigned(integer(my_cos(211)),16);
when x"0d4" => lut_sig <= to_unsigned(integer(my_cos(212)),16);
when x"0d5" => lut_sig <= to_unsigned(integer(my_cos(213)),16);
when x"0d6" => lut_sig <= to_unsigned(integer(my_cos(214)),16);
when x"0d7" => lut_sig <= to_unsigned(integer(my_cos(215)),16);
when x"0d8" => lut_sig <= to_unsigned(integer(my_cos(216)),16);
when x"0d9" => lut_sig <= to_unsigned(integer(my_cos(217)),16);
when x"0da" => lut_sig <= to_unsigned(integer(my_cos(218)),16);
when x"0db" => lut_sig <= to_unsigned(integer(my_cos(219)),16);
when x"0dc" => lut_sig <= to_unsigned(integer(my_cos(220)),16);
when x"0dd" => lut_sig <= to_unsigned(integer(my_cos(221)),16);
when x"0de" => lut_sig <= to_unsigned(integer(my_cos(222)),16);
when x"0df" => lut_sig <= to_unsigned(integer(my_cos(223)),16);
when x"0e0" => lut_sig <= to_unsigned(integer(my_cos(224)),16);
when x"0e1" => lut_sig <= to_unsigned(integer(my_cos(225)),16);
when x"0e2" => lut_sig <= to_unsigned(integer(my_cos(226)),16);
when x"0e3" => lut_sig <= to_unsigned(integer(my_cos(227)),16);
when x"0e4" => lut_sig <= to_unsigned(integer(my_cos(228)),16);
when x"0e5" => lut_sig <= to_unsigned(integer(my_cos(229)),16);
when x"0e6" => lut_sig <= to_unsigned(integer(my_cos(230)),16);
when x"0e7" => lut_sig <= to_unsigned(integer(my_cos(231)),16);
when x"0e8" => lut_sig <= to_unsigned(integer(my_cos(232)),16);
when x"0e9" => lut_sig <= to_unsigned(integer(my_cos(233)),16);
when x"0ea" => lut_sig <= to_unsigned(integer(my_cos(234)),16);
when x"0eb" => lut_sig <= to_unsigned(integer(my_cos(235)),16);
when x"0ec" => lut_sig <= to_unsigned(integer(my_cos(236)),16);
when x"0ed" => lut_sig <= to_unsigned(integer(my_cos(237)),16);
when x"0ee" => lut_sig <= to_unsigned(integer(my_cos(238)),16);
when x"0ef" => lut_sig <= to_unsigned(integer(my_cos(239)),16);
when x"0f0" => lut_sig <= to_unsigned(integer(my_cos(240)),16);
when x"0f1" => lut_sig <= to_unsigned(integer(my_cos(241)),16);
when x"0f2" => lut_sig <= to_unsigned(integer(my_cos(242)),16);
when x"0f3" => lut_sig <= to_unsigned(integer(my_cos(243)),16);
when x"0f4" => lut_sig <= to_unsigned(integer(my_cos(244)),16);
when x"0f5" => lut_sig <= to_unsigned(integer(my_cos(245)),16);
when x"0f6" => lut_sig <= to_unsigned(integer(my_cos(246)),16);
when x"0f7" => lut_sig <= to_unsigned(integer(my_cos(247)),16);
when x"0f8" => lut_sig <= to_unsigned(integer(my_cos(248)),16);
when x"0f9" => lut_sig <= to_unsigned(integer(my_cos(249)),16);
when x"0fa" => lut_sig <= to_unsigned(integer(my_cos(250)),16);
when x"0fb" => lut_sig <= to_unsigned(integer(my_cos(251)),16);
when x"0fc" => lut_sig <= to_unsigned(integer(my_cos(252)),16);
when x"0fd" => lut_sig <= to_unsigned(integer(my_cos(253)),16);
when x"0fe" => lut_sig <= to_unsigned(integer(my_cos(254)),16);
when x"0ff" => lut_sig <= to_unsigned(integer(my_cos(255)),16);
when x"100" => lut_sig <= to_unsigned(integer(my_cos(256)),16);
when x"101" => lut_sig <= to_unsigned(integer(my_cos(257)),16);
when x"102" => lut_sig <= to_unsigned(integer(my_cos(258)),16);
when x"103" => lut_sig <= to_unsigned(integer(my_cos(259)),16);
when x"104" => lut_sig <= to_unsigned(integer(my_cos(260)),16);
when x"105" => lut_sig <= to_unsigned(integer(my_cos(261)),16);
when x"106" => lut_sig <= to_unsigned(integer(my_cos(262)),16);
when x"107" => lut_sig <= to_unsigned(integer(my_cos(263)),16);
when x"108" => lut_sig <= to_unsigned(integer(my_cos(264)),16);
when x"109" => lut_sig <= to_unsigned(integer(my_cos(265)),16);
when x"10a" => lut_sig <= to_unsigned(integer(my_cos(266)),16);
when x"10b" => lut_sig <= to_unsigned(integer(my_cos(267)),16);
when x"10c" => lut_sig <= to_unsigned(integer(my_cos(268)),16);
when x"10d" => lut_sig <= to_unsigned(integer(my_cos(269)),16);
when x"10e" => lut_sig <= to_unsigned(integer(my_cos(270)),16);
when x"10f" => lut_sig <= to_unsigned(integer(my_cos(271)),16);
when x"110" => lut_sig <= to_unsigned(integer(my_cos(272)),16);
when x"111" => lut_sig <= to_unsigned(integer(my_cos(273)),16);
when x"112" => lut_sig <= to_unsigned(integer(my_cos(274)),16);
when x"113" => lut_sig <= to_unsigned(integer(my_cos(275)),16);
when x"114" => lut_sig <= to_unsigned(integer(my_cos(276)),16);
when x"115" => lut_sig <= to_unsigned(integer(my_cos(277)),16);
when x"116" => lut_sig <= to_unsigned(integer(my_cos(278)),16);
when x"117" => lut_sig <= to_unsigned(integer(my_cos(279)),16);
when x"118" => lut_sig <= to_unsigned(integer(my_cos(280)),16);
when x"119" => lut_sig <= to_unsigned(integer(my_cos(281)),16);
when x"11a" => lut_sig <= to_unsigned(integer(my_cos(282)),16);
when x"11b" => lut_sig <= to_unsigned(integer(my_cos(283)),16);
when x"11c" => lut_sig <= to_unsigned(integer(my_cos(284)),16);
when x"11d" => lut_sig <= to_unsigned(integer(my_cos(285)),16);
when x"11e" => lut_sig <= to_unsigned(integer(my_cos(286)),16);
when x"11f" => lut_sig <= to_unsigned(integer(my_cos(287)),16);
when x"120" => lut_sig <= to_unsigned(integer(my_cos(288)),16);
when x"121" => lut_sig <= to_unsigned(integer(my_cos(289)),16);
when x"122" => lut_sig <= to_unsigned(integer(my_cos(290)),16);
when x"123" => lut_sig <= to_unsigned(integer(my_cos(291)),16);
when x"124" => lut_sig <= to_unsigned(integer(my_cos(292)),16);
when x"125" => lut_sig <= to_unsigned(integer(my_cos(293)),16);
when x"126" => lut_sig <= to_unsigned(integer(my_cos(294)),16);
when x"127" => lut_sig <= to_unsigned(integer(my_cos(295)),16);
when x"128" => lut_sig <= to_unsigned(integer(my_cos(296)),16);
when x"129" => lut_sig <= to_unsigned(integer(my_cos(297)),16);
when x"12a" => lut_sig <= to_unsigned(integer(my_cos(298)),16);
when x"12b" => lut_sig <= to_unsigned(integer(my_cos(299)),16);
when x"12c" => lut_sig <= to_unsigned(integer(my_cos(300)),16);
when x"12d" => lut_sig <= to_unsigned(integer(my_cos(301)),16);
when x"12e" => lut_sig <= to_unsigned(integer(my_cos(302)),16);
when x"12f" => lut_sig <= to_unsigned(integer(my_cos(303)),16);
when x"130" => lut_sig <= to_unsigned(integer(my_cos(304)),16);
when x"131" => lut_sig <= to_unsigned(integer(my_cos(305)),16);
when x"132" => lut_sig <= to_unsigned(integer(my_cos(306)),16);
when x"133" => lut_sig <= to_unsigned(integer(my_cos(307)),16);
when x"134" => lut_sig <= to_unsigned(integer(my_cos(308)),16);
when x"135" => lut_sig <= to_unsigned(integer(my_cos(309)),16);
when x"136" => lut_sig <= to_unsigned(integer(my_cos(310)),16);
when x"137" => lut_sig <= to_unsigned(integer(my_cos(311)),16);
when x"138" => lut_sig <= to_unsigned(integer(my_cos(312)),16);
when x"139" => lut_sig <= to_unsigned(integer(my_cos(313)),16);
when x"13a" => lut_sig <= to_unsigned(integer(my_cos(314)),16);
when x"13b" => lut_sig <= to_unsigned(integer(my_cos(315)),16);
when x"13c" => lut_sig <= to_unsigned(integer(my_cos(316)),16);
when x"13d" => lut_sig <= to_unsigned(integer(my_cos(317)),16);
when x"13e" => lut_sig <= to_unsigned(integer(my_cos(318)),16);
when x"13f" => lut_sig <= to_unsigned(integer(my_cos(319)),16);
when x"140" => lut_sig <= to_unsigned(integer(my_cos(320)),16);
when x"141" => lut_sig <= to_unsigned(integer(my_cos(321)),16);
when x"142" => lut_sig <= to_unsigned(integer(my_cos(322)),16);
when x"143" => lut_sig <= to_unsigned(integer(my_cos(323)),16);
when x"144" => lut_sig <= to_unsigned(integer(my_cos(324)),16);
when x"145" => lut_sig <= to_unsigned(integer(my_cos(325)),16);
when x"146" => lut_sig <= to_unsigned(integer(my_cos(326)),16);
when x"147" => lut_sig <= to_unsigned(integer(my_cos(327)),16);
when x"148" => lut_sig <= to_unsigned(integer(my_cos(328)),16);
when x"149" => lut_sig <= to_unsigned(integer(my_cos(329)),16);
when x"14a" => lut_sig <= to_unsigned(integer(my_cos(330)),16);
when x"14b" => lut_sig <= to_unsigned(integer(my_cos(331)),16);
when x"14c" => lut_sig <= to_unsigned(integer(my_cos(332)),16);
when x"14d" => lut_sig <= to_unsigned(integer(my_cos(333)),16);
when x"14e" => lut_sig <= to_unsigned(integer(my_cos(334)),16);
when x"14f" => lut_sig <= to_unsigned(integer(my_cos(335)),16);
when x"150" => lut_sig <= to_unsigned(integer(my_cos(336)),16);
when x"151" => lut_sig <= to_unsigned(integer(my_cos(337)),16);
when x"152" => lut_sig <= to_unsigned(integer(my_cos(338)),16);
when x"153" => lut_sig <= to_unsigned(integer(my_cos(339)),16);
when x"154" => lut_sig <= to_unsigned(integer(my_cos(340)),16);
when x"155" => lut_sig <= to_unsigned(integer(my_cos(341)),16);
when x"156" => lut_sig <= to_unsigned(integer(my_cos(342)),16);
when x"157" => lut_sig <= to_unsigned(integer(my_cos(343)),16);
when x"158" => lut_sig <= to_unsigned(integer(my_cos(344)),16);
when x"159" => lut_sig <= to_unsigned(integer(my_cos(345)),16);
when x"15a" => lut_sig <= to_unsigned(integer(my_cos(346)),16);
when x"15b" => lut_sig <= to_unsigned(integer(my_cos(347)),16);
when x"15c" => lut_sig <= to_unsigned(integer(my_cos(348)),16);
when x"15d" => lut_sig <= to_unsigned(integer(my_cos(349)),16);
when x"15e" => lut_sig <= to_unsigned(integer(my_cos(350)),16);
when x"15f" => lut_sig <= to_unsigned(integer(my_cos(351)),16);
when x"160" => lut_sig <= to_unsigned(integer(my_cos(352)),16);
when x"161" => lut_sig <= to_unsigned(integer(my_cos(353)),16);
when x"162" => lut_sig <= to_unsigned(integer(my_cos(354)),16);
when x"163" => lut_sig <= to_unsigned(integer(my_cos(355)),16);
when x"164" => lut_sig <= to_unsigned(integer(my_cos(356)),16);
when x"165" => lut_sig <= to_unsigned(integer(my_cos(357)),16);
when x"166" => lut_sig <= to_unsigned(integer(my_cos(358)),16);
when x"167" => lut_sig <= to_unsigned(integer(my_cos(359)),16);
when x"168" => lut_sig <= to_unsigned(integer(my_cos(360)),16);
when x"169" => lut_sig <= to_unsigned(integer(my_cos(361)),16);
when x"16a" => lut_sig <= to_unsigned(integer(my_cos(362)),16);
when x"16b" => lut_sig <= to_unsigned(integer(my_cos(363)),16);
when x"16c" => lut_sig <= to_unsigned(integer(my_cos(364)),16);
when x"16d" => lut_sig <= to_unsigned(integer(my_cos(365)),16);
when x"16e" => lut_sig <= to_unsigned(integer(my_cos(366)),16);
when x"16f" => lut_sig <= to_unsigned(integer(my_cos(367)),16);
when x"170" => lut_sig <= to_unsigned(integer(my_cos(368)),16);
when x"171" => lut_sig <= to_unsigned(integer(my_cos(369)),16);
when x"172" => lut_sig <= to_unsigned(integer(my_cos(370)),16);
when x"173" => lut_sig <= to_unsigned(integer(my_cos(371)),16);
when x"174" => lut_sig <= to_unsigned(integer(my_cos(372)),16);
when x"175" => lut_sig <= to_unsigned(integer(my_cos(373)),16);
when x"176" => lut_sig <= to_unsigned(integer(my_cos(374)),16);
when x"177" => lut_sig <= to_unsigned(integer(my_cos(375)),16);
when x"178" => lut_sig <= to_unsigned(integer(my_cos(376)),16);
when x"179" => lut_sig <= to_unsigned(integer(my_cos(377)),16);
when x"17a" => lut_sig <= to_unsigned(integer(my_cos(378)),16);
when x"17b" => lut_sig <= to_unsigned(integer(my_cos(379)),16);
when x"17c" => lut_sig <= to_unsigned(integer(my_cos(380)),16);
when x"17d" => lut_sig <= to_unsigned(integer(my_cos(381)),16);
when x"17e" => lut_sig <= to_unsigned(integer(my_cos(382)),16);
when x"17f" => lut_sig <= to_unsigned(integer(my_cos(383)),16);
when x"180" => lut_sig <= to_unsigned(integer(my_cos(384)),16);
when x"181" => lut_sig <= to_unsigned(integer(my_cos(385)),16);
when x"182" => lut_sig <= to_unsigned(integer(my_cos(386)),16);
when x"183" => lut_sig <= to_unsigned(integer(my_cos(387)),16);
when x"184" => lut_sig <= to_unsigned(integer(my_cos(388)),16);
when x"185" => lut_sig <= to_unsigned(integer(my_cos(389)),16);
when x"186" => lut_sig <= to_unsigned(integer(my_cos(390)),16);
when x"187" => lut_sig <= to_unsigned(integer(my_cos(391)),16);
when x"188" => lut_sig <= to_unsigned(integer(my_cos(392)),16);
when x"189" => lut_sig <= to_unsigned(integer(my_cos(393)),16);
when x"18a" => lut_sig <= to_unsigned(integer(my_cos(394)),16);
when x"18b" => lut_sig <= to_unsigned(integer(my_cos(395)),16);
when x"18c" => lut_sig <= to_unsigned(integer(my_cos(396)),16);
when x"18d" => lut_sig <= to_unsigned(integer(my_cos(397)),16);
when x"18e" => lut_sig <= to_unsigned(integer(my_cos(398)),16);
when x"18f" => lut_sig <= to_unsigned(integer(my_cos(399)),16);
when x"190" => lut_sig <= to_unsigned(integer(my_cos(400)),16);
when x"191" => lut_sig <= to_unsigned(integer(my_cos(401)),16);
when x"192" => lut_sig <= to_unsigned(integer(my_cos(402)),16);
when x"193" => lut_sig <= to_unsigned(integer(my_cos(403)),16);
when x"194" => lut_sig <= to_unsigned(integer(my_cos(404)),16);
when x"195" => lut_sig <= to_unsigned(integer(my_cos(405)),16);
when x"196" => lut_sig <= to_unsigned(integer(my_cos(406)),16);
when x"197" => lut_sig <= to_unsigned(integer(my_cos(407)),16);
when x"198" => lut_sig <= to_unsigned(integer(my_cos(408)),16);
when x"199" => lut_sig <= to_unsigned(integer(my_cos(409)),16);
when x"19a" => lut_sig <= to_unsigned(integer(my_cos(410)),16);
when x"19b" => lut_sig <= to_unsigned(integer(my_cos(411)),16);
when x"19c" => lut_sig <= to_unsigned(integer(my_cos(412)),16);
when x"19d" => lut_sig <= to_unsigned(integer(my_cos(413)),16);
when x"19e" => lut_sig <= to_unsigned(integer(my_cos(414)),16);
when x"19f" => lut_sig <= to_unsigned(integer(my_cos(415)),16);
when x"1a0" => lut_sig <= to_unsigned(integer(my_cos(416)),16);
when x"1a1" => lut_sig <= to_unsigned(integer(my_cos(417)),16);
when x"1a2" => lut_sig <= to_unsigned(integer(my_cos(418)),16);
when x"1a3" => lut_sig <= to_unsigned(integer(my_cos(419)),16);
when x"1a4" => lut_sig <= to_unsigned(integer(my_cos(420)),16);
when x"1a5" => lut_sig <= to_unsigned(integer(my_cos(421)),16);
when x"1a6" => lut_sig <= to_unsigned(integer(my_cos(422)),16);
when x"1a7" => lut_sig <= to_unsigned(integer(my_cos(423)),16);
when x"1a8" => lut_sig <= to_unsigned(integer(my_cos(424)),16);
when x"1a9" => lut_sig <= to_unsigned(integer(my_cos(425)),16);
when x"1aa" => lut_sig <= to_unsigned(integer(my_cos(426)),16);
when x"1ab" => lut_sig <= to_unsigned(integer(my_cos(427)),16);
when x"1ac" => lut_sig <= to_unsigned(integer(my_cos(428)),16);
when x"1ad" => lut_sig <= to_unsigned(integer(my_cos(429)),16);
when x"1ae" => lut_sig <= to_unsigned(integer(my_cos(430)),16);
when x"1af" => lut_sig <= to_unsigned(integer(my_cos(431)),16);
when x"1b0" => lut_sig <= to_unsigned(integer(my_cos(432)),16);
when x"1b1" => lut_sig <= to_unsigned(integer(my_cos(433)),16);
when x"1b2" => lut_sig <= to_unsigned(integer(my_cos(434)),16);
when x"1b3" => lut_sig <= to_unsigned(integer(my_cos(435)),16);
when x"1b4" => lut_sig <= to_unsigned(integer(my_cos(436)),16);
when x"1b5" => lut_sig <= to_unsigned(integer(my_cos(437)),16);
when x"1b6" => lut_sig <= to_unsigned(integer(my_cos(438)),16);
when x"1b7" => lut_sig <= to_unsigned(integer(my_cos(439)),16);
when x"1b8" => lut_sig <= to_unsigned(integer(my_cos(440)),16);
when x"1b9" => lut_sig <= to_unsigned(integer(my_cos(441)),16);
when x"1ba" => lut_sig <= to_unsigned(integer(my_cos(442)),16);
when x"1bb" => lut_sig <= to_unsigned(integer(my_cos(443)),16);
when x"1bc" => lut_sig <= to_unsigned(integer(my_cos(444)),16);
when x"1bd" => lut_sig <= to_unsigned(integer(my_cos(445)),16);
when x"1be" => lut_sig <= to_unsigned(integer(my_cos(446)),16);
when x"1bf" => lut_sig <= to_unsigned(integer(my_cos(447)),16);
when x"1c0" => lut_sig <= to_unsigned(integer(my_cos(448)),16);
when x"1c1" => lut_sig <= to_unsigned(integer(my_cos(449)),16);
when x"1c2" => lut_sig <= to_unsigned(integer(my_cos(450)),16);
when x"1c3" => lut_sig <= to_unsigned(integer(my_cos(451)),16);
when x"1c4" => lut_sig <= to_unsigned(integer(my_cos(452)),16);
when x"1c5" => lut_sig <= to_unsigned(integer(my_cos(453)),16);
when x"1c6" => lut_sig <= to_unsigned(integer(my_cos(454)),16);
when x"1c7" => lut_sig <= to_unsigned(integer(my_cos(455)),16);
when x"1c8" => lut_sig <= to_unsigned(integer(my_cos(456)),16);
when x"1c9" => lut_sig <= to_unsigned(integer(my_cos(457)),16);
when x"1ca" => lut_sig <= to_unsigned(integer(my_cos(458)),16);
when x"1cb" => lut_sig <= to_unsigned(integer(my_cos(459)),16);
when x"1cc" => lut_sig <= to_unsigned(integer(my_cos(460)),16);
when x"1cd" => lut_sig <= to_unsigned(integer(my_cos(461)),16);
when x"1ce" => lut_sig <= to_unsigned(integer(my_cos(462)),16);
when x"1cf" => lut_sig <= to_unsigned(integer(my_cos(463)),16);
when x"1d0" => lut_sig <= to_unsigned(integer(my_cos(464)),16);
when x"1d1" => lut_sig <= to_unsigned(integer(my_cos(465)),16);
when x"1d2" => lut_sig <= to_unsigned(integer(my_cos(466)),16);
when x"1d3" => lut_sig <= to_unsigned(integer(my_cos(467)),16);
when x"1d4" => lut_sig <= to_unsigned(integer(my_cos(468)),16);
when x"1d5" => lut_sig <= to_unsigned(integer(my_cos(469)),16);
when x"1d6" => lut_sig <= to_unsigned(integer(my_cos(470)),16);
when x"1d7" => lut_sig <= to_unsigned(integer(my_cos(471)),16);
when x"1d8" => lut_sig <= to_unsigned(integer(my_cos(472)),16);
when x"1d9" => lut_sig <= to_unsigned(integer(my_cos(473)),16);
when x"1da" => lut_sig <= to_unsigned(integer(my_cos(474)),16);
when x"1db" => lut_sig <= to_unsigned(integer(my_cos(475)),16);
when x"1dc" => lut_sig <= to_unsigned(integer(my_cos(476)),16);
when x"1dd" => lut_sig <= to_unsigned(integer(my_cos(477)),16);
when x"1de" => lut_sig <= to_unsigned(integer(my_cos(478)),16);
when x"1df" => lut_sig <= to_unsigned(integer(my_cos(479)),16);
when x"1e0" => lut_sig <= to_unsigned(integer(my_cos(480)),16);
when x"1e1" => lut_sig <= to_unsigned(integer(my_cos(481)),16);
when x"1e2" => lut_sig <= to_unsigned(integer(my_cos(482)),16);
when x"1e3" => lut_sig <= to_unsigned(integer(my_cos(483)),16);
when x"1e4" => lut_sig <= to_unsigned(integer(my_cos(484)),16);
when x"1e5" => lut_sig <= to_unsigned(integer(my_cos(485)),16);
when x"1e6" => lut_sig <= to_unsigned(integer(my_cos(486)),16);
when x"1e7" => lut_sig <= to_unsigned(integer(my_cos(487)),16);
when x"1e8" => lut_sig <= to_unsigned(integer(my_cos(488)),16);
when x"1e9" => lut_sig <= to_unsigned(integer(my_cos(489)),16);
when x"1ea" => lut_sig <= to_unsigned(integer(my_cos(490)),16);
when x"1eb" => lut_sig <= to_unsigned(integer(my_cos(491)),16);
when x"1ec" => lut_sig <= to_unsigned(integer(my_cos(492)),16);
when x"1ed" => lut_sig <= to_unsigned(integer(my_cos(493)),16);
when x"1ee" => lut_sig <= to_unsigned(integer(my_cos(494)),16);
when x"1ef" => lut_sig <= to_unsigned(integer(my_cos(495)),16);
when x"1f0" => lut_sig <= to_unsigned(integer(my_cos(496)),16);
when x"1f1" => lut_sig <= to_unsigned(integer(my_cos(497)),16);
when x"1f2" => lut_sig <= to_unsigned(integer(my_cos(498)),16);
when x"1f3" => lut_sig <= to_unsigned(integer(my_cos(499)),16);
when x"1f4" => lut_sig <= to_unsigned(integer(my_cos(500)),16);
when x"1f5" => lut_sig <= to_unsigned(integer(my_cos(501)),16);
when x"1f6" => lut_sig <= to_unsigned(integer(my_cos(502)),16);
when x"1f7" => lut_sig <= to_unsigned(integer(my_cos(503)),16);
when x"1f8" => lut_sig <= to_unsigned(integer(my_cos(504)),16);
when x"1f9" => lut_sig <= to_unsigned(integer(my_cos(505)),16);
when x"1fa" => lut_sig <= to_unsigned(integer(my_cos(506)),16);
when x"1fb" => lut_sig <= to_unsigned(integer(my_cos(507)),16);
when x"1fc" => lut_sig <= to_unsigned(integer(my_cos(508)),16);
when x"1fd" => lut_sig <= to_unsigned(integer(my_cos(509)),16);
when x"1fe" => lut_sig <= to_unsigned(integer(my_cos(510)),16);
when x"1ff" => lut_sig <= to_unsigned(integer(my_cos(511)),16);
when x"200" => lut_sig <= to_unsigned(integer(my_cos(512)),16);
when x"201" => lut_sig <= to_unsigned(integer(my_cos(513)),16);
when x"202" => lut_sig <= to_unsigned(integer(my_cos(514)),16);
when x"203" => lut_sig <= to_unsigned(integer(my_cos(515)),16);
when x"204" => lut_sig <= to_unsigned(integer(my_cos(516)),16);
when x"205" => lut_sig <= to_unsigned(integer(my_cos(517)),16);
when x"206" => lut_sig <= to_unsigned(integer(my_cos(518)),16);
when x"207" => lut_sig <= to_unsigned(integer(my_cos(519)),16);
when x"208" => lut_sig <= to_unsigned(integer(my_cos(520)),16);
when x"209" => lut_sig <= to_unsigned(integer(my_cos(521)),16);
when x"20a" => lut_sig <= to_unsigned(integer(my_cos(522)),16);
when x"20b" => lut_sig <= to_unsigned(integer(my_cos(523)),16);
when x"20c" => lut_sig <= to_unsigned(integer(my_cos(524)),16);
when x"20d" => lut_sig <= to_unsigned(integer(my_cos(525)),16);
when x"20e" => lut_sig <= to_unsigned(integer(my_cos(526)),16);
when x"20f" => lut_sig <= to_unsigned(integer(my_cos(527)),16);
when x"210" => lut_sig <= to_unsigned(integer(my_cos(528)),16);
when x"211" => lut_sig <= to_unsigned(integer(my_cos(529)),16);
when x"212" => lut_sig <= to_unsigned(integer(my_cos(530)),16);
when x"213" => lut_sig <= to_unsigned(integer(my_cos(531)),16);
when x"214" => lut_sig <= to_unsigned(integer(my_cos(532)),16);
when x"215" => lut_sig <= to_unsigned(integer(my_cos(533)),16);
when x"216" => lut_sig <= to_unsigned(integer(my_cos(534)),16);
when x"217" => lut_sig <= to_unsigned(integer(my_cos(535)),16);
when x"218" => lut_sig <= to_unsigned(integer(my_cos(536)),16);
when x"219" => lut_sig <= to_unsigned(integer(my_cos(537)),16);
when x"21a" => lut_sig <= to_unsigned(integer(my_cos(538)),16);
when x"21b" => lut_sig <= to_unsigned(integer(my_cos(539)),16);
when x"21c" => lut_sig <= to_unsigned(integer(my_cos(540)),16);
when x"21d" => lut_sig <= to_unsigned(integer(my_cos(541)),16);
when x"21e" => lut_sig <= to_unsigned(integer(my_cos(542)),16);
when x"21f" => lut_sig <= to_unsigned(integer(my_cos(543)),16);
when x"220" => lut_sig <= to_unsigned(integer(my_cos(544)),16);
when x"221" => lut_sig <= to_unsigned(integer(my_cos(545)),16);
when x"222" => lut_sig <= to_unsigned(integer(my_cos(546)),16);
when x"223" => lut_sig <= to_unsigned(integer(my_cos(547)),16);
when x"224" => lut_sig <= to_unsigned(integer(my_cos(548)),16);
when x"225" => lut_sig <= to_unsigned(integer(my_cos(549)),16);
when x"226" => lut_sig <= to_unsigned(integer(my_cos(550)),16);
when x"227" => lut_sig <= to_unsigned(integer(my_cos(551)),16);
when x"228" => lut_sig <= to_unsigned(integer(my_cos(552)),16);
when x"229" => lut_sig <= to_unsigned(integer(my_cos(553)),16);
when x"22a" => lut_sig <= to_unsigned(integer(my_cos(554)),16);
when x"22b" => lut_sig <= to_unsigned(integer(my_cos(555)),16);
when x"22c" => lut_sig <= to_unsigned(integer(my_cos(556)),16);
when x"22d" => lut_sig <= to_unsigned(integer(my_cos(557)),16);
when x"22e" => lut_sig <= to_unsigned(integer(my_cos(558)),16);
when x"22f" => lut_sig <= to_unsigned(integer(my_cos(559)),16);
when x"230" => lut_sig <= to_unsigned(integer(my_cos(560)),16);
when x"231" => lut_sig <= to_unsigned(integer(my_cos(561)),16);
when x"232" => lut_sig <= to_unsigned(integer(my_cos(562)),16);
when x"233" => lut_sig <= to_unsigned(integer(my_cos(563)),16);
when x"234" => lut_sig <= to_unsigned(integer(my_cos(564)),16);
when x"235" => lut_sig <= to_unsigned(integer(my_cos(565)),16);
when x"236" => lut_sig <= to_unsigned(integer(my_cos(566)),16);
when x"237" => lut_sig <= to_unsigned(integer(my_cos(567)),16);
when x"238" => lut_sig <= to_unsigned(integer(my_cos(568)),16);
when x"239" => lut_sig <= to_unsigned(integer(my_cos(569)),16);
when x"23a" => lut_sig <= to_unsigned(integer(my_cos(570)),16);
when x"23b" => lut_sig <= to_unsigned(integer(my_cos(571)),16);
when x"23c" => lut_sig <= to_unsigned(integer(my_cos(572)),16);
when x"23d" => lut_sig <= to_unsigned(integer(my_cos(573)),16);
when x"23e" => lut_sig <= to_unsigned(integer(my_cos(574)),16);
when x"23f" => lut_sig <= to_unsigned(integer(my_cos(575)),16);
when x"240" => lut_sig <= to_unsigned(integer(my_cos(576)),16);
when x"241" => lut_sig <= to_unsigned(integer(my_cos(577)),16);
when x"242" => lut_sig <= to_unsigned(integer(my_cos(578)),16);
when x"243" => lut_sig <= to_unsigned(integer(my_cos(579)),16);
when x"244" => lut_sig <= to_unsigned(integer(my_cos(580)),16);
when x"245" => lut_sig <= to_unsigned(integer(my_cos(581)),16);
when x"246" => lut_sig <= to_unsigned(integer(my_cos(582)),16);
when x"247" => lut_sig <= to_unsigned(integer(my_cos(583)),16);
when x"248" => lut_sig <= to_unsigned(integer(my_cos(584)),16);
when x"249" => lut_sig <= to_unsigned(integer(my_cos(585)),16);
when x"24a" => lut_sig <= to_unsigned(integer(my_cos(586)),16);
when x"24b" => lut_sig <= to_unsigned(integer(my_cos(587)),16);
when x"24c" => lut_sig <= to_unsigned(integer(my_cos(588)),16);
when x"24d" => lut_sig <= to_unsigned(integer(my_cos(589)),16);
when x"24e" => lut_sig <= to_unsigned(integer(my_cos(590)),16);
when x"24f" => lut_sig <= to_unsigned(integer(my_cos(591)),16);
when x"250" => lut_sig <= to_unsigned(integer(my_cos(592)),16);
when x"251" => lut_sig <= to_unsigned(integer(my_cos(593)),16);
when x"252" => lut_sig <= to_unsigned(integer(my_cos(594)),16);
when x"253" => lut_sig <= to_unsigned(integer(my_cos(595)),16);
when x"254" => lut_sig <= to_unsigned(integer(my_cos(596)),16);
when x"255" => lut_sig <= to_unsigned(integer(my_cos(597)),16);
when x"256" => lut_sig <= to_unsigned(integer(my_cos(598)),16);
when x"257" => lut_sig <= to_unsigned(integer(my_cos(599)),16);
when x"258" => lut_sig <= to_unsigned(integer(my_cos(600)),16);
when x"259" => lut_sig <= to_unsigned(integer(my_cos(601)),16);
when x"25a" => lut_sig <= to_unsigned(integer(my_cos(602)),16);
when x"25b" => lut_sig <= to_unsigned(integer(my_cos(603)),16);
when x"25c" => lut_sig <= to_unsigned(integer(my_cos(604)),16);
when x"25d" => lut_sig <= to_unsigned(integer(my_cos(605)),16);
when x"25e" => lut_sig <= to_unsigned(integer(my_cos(606)),16);
when x"25f" => lut_sig <= to_unsigned(integer(my_cos(607)),16);
when x"260" => lut_sig <= to_unsigned(integer(my_cos(608)),16);
when x"261" => lut_sig <= to_unsigned(integer(my_cos(609)),16);
when x"262" => lut_sig <= to_unsigned(integer(my_cos(610)),16);
when x"263" => lut_sig <= to_unsigned(integer(my_cos(611)),16);
when x"264" => lut_sig <= to_unsigned(integer(my_cos(612)),16);
when x"265" => lut_sig <= to_unsigned(integer(my_cos(613)),16);
when x"266" => lut_sig <= to_unsigned(integer(my_cos(614)),16);
when x"267" => lut_sig <= to_unsigned(integer(my_cos(615)),16);
when x"268" => lut_sig <= to_unsigned(integer(my_cos(616)),16);
when x"269" => lut_sig <= to_unsigned(integer(my_cos(617)),16);
when x"26a" => lut_sig <= to_unsigned(integer(my_cos(618)),16);
when x"26b" => lut_sig <= to_unsigned(integer(my_cos(619)),16);
when x"26c" => lut_sig <= to_unsigned(integer(my_cos(620)),16);
when x"26d" => lut_sig <= to_unsigned(integer(my_cos(621)),16);
when x"26e" => lut_sig <= to_unsigned(integer(my_cos(622)),16);
when x"26f" => lut_sig <= to_unsigned(integer(my_cos(623)),16);
when x"270" => lut_sig <= to_unsigned(integer(my_cos(624)),16);
when x"271" => lut_sig <= to_unsigned(integer(my_cos(625)),16);
when x"272" => lut_sig <= to_unsigned(integer(my_cos(626)),16);
when x"273" => lut_sig <= to_unsigned(integer(my_cos(627)),16);
when x"274" => lut_sig <= to_unsigned(integer(my_cos(628)),16);
when x"275" => lut_sig <= to_unsigned(integer(my_cos(629)),16);
when x"276" => lut_sig <= to_unsigned(integer(my_cos(630)),16);
when x"277" => lut_sig <= to_unsigned(integer(my_cos(631)),16);
when x"278" => lut_sig <= to_unsigned(integer(my_cos(632)),16);
when x"279" => lut_sig <= to_unsigned(integer(my_cos(633)),16);
when x"27a" => lut_sig <= to_unsigned(integer(my_cos(634)),16);
when x"27b" => lut_sig <= to_unsigned(integer(my_cos(635)),16);
when x"27c" => lut_sig <= to_unsigned(integer(my_cos(636)),16);
when x"27d" => lut_sig <= to_unsigned(integer(my_cos(637)),16);
when x"27e" => lut_sig <= to_unsigned(integer(my_cos(638)),16);
when x"27f" => lut_sig <= to_unsigned(integer(my_cos(639)),16);
when x"280" => lut_sig <= to_unsigned(integer(my_cos(640)),16);
when x"281" => lut_sig <= to_unsigned(integer(my_cos(641)),16);
when x"282" => lut_sig <= to_unsigned(integer(my_cos(642)),16);
when x"283" => lut_sig <= to_unsigned(integer(my_cos(643)),16);
when x"284" => lut_sig <= to_unsigned(integer(my_cos(644)),16);
when x"285" => lut_sig <= to_unsigned(integer(my_cos(645)),16);
when x"286" => lut_sig <= to_unsigned(integer(my_cos(646)),16);
when x"287" => lut_sig <= to_unsigned(integer(my_cos(647)),16);
when x"288" => lut_sig <= to_unsigned(integer(my_cos(648)),16);
when x"289" => lut_sig <= to_unsigned(integer(my_cos(649)),16);
when x"28a" => lut_sig <= to_unsigned(integer(my_cos(650)),16);
when x"28b" => lut_sig <= to_unsigned(integer(my_cos(651)),16);
when x"28c" => lut_sig <= to_unsigned(integer(my_cos(652)),16);
when x"28d" => lut_sig <= to_unsigned(integer(my_cos(653)),16);
when x"28e" => lut_sig <= to_unsigned(integer(my_cos(654)),16);
when x"28f" => lut_sig <= to_unsigned(integer(my_cos(655)),16);
when x"290" => lut_sig <= to_unsigned(integer(my_cos(656)),16);
when x"291" => lut_sig <= to_unsigned(integer(my_cos(657)),16);
when x"292" => lut_sig <= to_unsigned(integer(my_cos(658)),16);
when x"293" => lut_sig <= to_unsigned(integer(my_cos(659)),16);
when x"294" => lut_sig <= to_unsigned(integer(my_cos(660)),16);
when x"295" => lut_sig <= to_unsigned(integer(my_cos(661)),16);
when x"296" => lut_sig <= to_unsigned(integer(my_cos(662)),16);
when x"297" => lut_sig <= to_unsigned(integer(my_cos(663)),16);
when x"298" => lut_sig <= to_unsigned(integer(my_cos(664)),16);
when x"299" => lut_sig <= to_unsigned(integer(my_cos(665)),16);
when x"29a" => lut_sig <= to_unsigned(integer(my_cos(666)),16);
when x"29b" => lut_sig <= to_unsigned(integer(my_cos(667)),16);
when x"29c" => lut_sig <= to_unsigned(integer(my_cos(668)),16);
when x"29d" => lut_sig <= to_unsigned(integer(my_cos(669)),16);
when x"29e" => lut_sig <= to_unsigned(integer(my_cos(670)),16);
when x"29f" => lut_sig <= to_unsigned(integer(my_cos(671)),16);
when x"2a0" => lut_sig <= to_unsigned(integer(my_cos(672)),16);
when x"2a1" => lut_sig <= to_unsigned(integer(my_cos(673)),16);
when x"2a2" => lut_sig <= to_unsigned(integer(my_cos(674)),16);
when x"2a3" => lut_sig <= to_unsigned(integer(my_cos(675)),16);
when x"2a4" => lut_sig <= to_unsigned(integer(my_cos(676)),16);
when x"2a5" => lut_sig <= to_unsigned(integer(my_cos(677)),16);
when x"2a6" => lut_sig <= to_unsigned(integer(my_cos(678)),16);
when x"2a7" => lut_sig <= to_unsigned(integer(my_cos(679)),16);
when x"2a8" => lut_sig <= to_unsigned(integer(my_cos(680)),16);
when x"2a9" => lut_sig <= to_unsigned(integer(my_cos(681)),16);
when x"2aa" => lut_sig <= to_unsigned(integer(my_cos(682)),16);
when x"2ab" => lut_sig <= to_unsigned(integer(my_cos(683)),16);
when x"2ac" => lut_sig <= to_unsigned(integer(my_cos(684)),16);
when x"2ad" => lut_sig <= to_unsigned(integer(my_cos(685)),16);
when x"2ae" => lut_sig <= to_unsigned(integer(my_cos(686)),16);
when x"2af" => lut_sig <= to_unsigned(integer(my_cos(687)),16);
when x"2b0" => lut_sig <= to_unsigned(integer(my_cos(688)),16);
when x"2b1" => lut_sig <= to_unsigned(integer(my_cos(689)),16);
when x"2b2" => lut_sig <= to_unsigned(integer(my_cos(690)),16);
when x"2b3" => lut_sig <= to_unsigned(integer(my_cos(691)),16);
when x"2b4" => lut_sig <= to_unsigned(integer(my_cos(692)),16);
when x"2b5" => lut_sig <= to_unsigned(integer(my_cos(693)),16);
when x"2b6" => lut_sig <= to_unsigned(integer(my_cos(694)),16);
when x"2b7" => lut_sig <= to_unsigned(integer(my_cos(695)),16);
when x"2b8" => lut_sig <= to_unsigned(integer(my_cos(696)),16);
when x"2b9" => lut_sig <= to_unsigned(integer(my_cos(697)),16);
when x"2ba" => lut_sig <= to_unsigned(integer(my_cos(698)),16);
when x"2bb" => lut_sig <= to_unsigned(integer(my_cos(699)),16);
when x"2bc" => lut_sig <= to_unsigned(integer(my_cos(700)),16);
when x"2bd" => lut_sig <= to_unsigned(integer(my_cos(701)),16);
when x"2be" => lut_sig <= to_unsigned(integer(my_cos(702)),16);
when x"2bf" => lut_sig <= to_unsigned(integer(my_cos(703)),16);
when x"2c0" => lut_sig <= to_unsigned(integer(my_cos(704)),16);
when x"2c1" => lut_sig <= to_unsigned(integer(my_cos(705)),16);
when x"2c2" => lut_sig <= to_unsigned(integer(my_cos(706)),16);
when x"2c3" => lut_sig <= to_unsigned(integer(my_cos(707)),16);
when x"2c4" => lut_sig <= to_unsigned(integer(my_cos(708)),16);
when x"2c5" => lut_sig <= to_unsigned(integer(my_cos(709)),16);
when x"2c6" => lut_sig <= to_unsigned(integer(my_cos(710)),16);
when x"2c7" => lut_sig <= to_unsigned(integer(my_cos(711)),16);
when x"2c8" => lut_sig <= to_unsigned(integer(my_cos(712)),16);
when x"2c9" => lut_sig <= to_unsigned(integer(my_cos(713)),16);
when x"2ca" => lut_sig <= to_unsigned(integer(my_cos(714)),16);
when x"2cb" => lut_sig <= to_unsigned(integer(my_cos(715)),16);
when x"2cc" => lut_sig <= to_unsigned(integer(my_cos(716)),16);
when x"2cd" => lut_sig <= to_unsigned(integer(my_cos(717)),16);
when x"2ce" => lut_sig <= to_unsigned(integer(my_cos(718)),16);
when x"2cf" => lut_sig <= to_unsigned(integer(my_cos(719)),16);
when x"2d0" => lut_sig <= to_unsigned(integer(my_cos(720)),16);
when x"2d1" => lut_sig <= to_unsigned(integer(my_cos(721)),16);
when x"2d2" => lut_sig <= to_unsigned(integer(my_cos(722)),16);
when x"2d3" => lut_sig <= to_unsigned(integer(my_cos(723)),16);
when x"2d4" => lut_sig <= to_unsigned(integer(my_cos(724)),16);
when x"2d5" => lut_sig <= to_unsigned(integer(my_cos(725)),16);
when x"2d6" => lut_sig <= to_unsigned(integer(my_cos(726)),16);
when x"2d7" => lut_sig <= to_unsigned(integer(my_cos(727)),16);
when x"2d8" => lut_sig <= to_unsigned(integer(my_cos(728)),16);
when x"2d9" => lut_sig <= to_unsigned(integer(my_cos(729)),16);
when x"2da" => lut_sig <= to_unsigned(integer(my_cos(730)),16);
when x"2db" => lut_sig <= to_unsigned(integer(my_cos(731)),16);
when x"2dc" => lut_sig <= to_unsigned(integer(my_cos(732)),16);
when x"2dd" => lut_sig <= to_unsigned(integer(my_cos(733)),16);
when x"2de" => lut_sig <= to_unsigned(integer(my_cos(734)),16);
when x"2df" => lut_sig <= to_unsigned(integer(my_cos(735)),16);
when x"2e0" => lut_sig <= to_unsigned(integer(my_cos(736)),16);
when x"2e1" => lut_sig <= to_unsigned(integer(my_cos(737)),16);
when x"2e2" => lut_sig <= to_unsigned(integer(my_cos(738)),16);
when x"2e3" => lut_sig <= to_unsigned(integer(my_cos(739)),16);
when x"2e4" => lut_sig <= to_unsigned(integer(my_cos(740)),16);
when x"2e5" => lut_sig <= to_unsigned(integer(my_cos(741)),16);
when x"2e6" => lut_sig <= to_unsigned(integer(my_cos(742)),16);
when x"2e7" => lut_sig <= to_unsigned(integer(my_cos(743)),16);
when x"2e8" => lut_sig <= to_unsigned(integer(my_cos(744)),16);
when x"2e9" => lut_sig <= to_unsigned(integer(my_cos(745)),16);
when x"2ea" => lut_sig <= to_unsigned(integer(my_cos(746)),16);
when x"2eb" => lut_sig <= to_unsigned(integer(my_cos(747)),16);
when x"2ec" => lut_sig <= to_unsigned(integer(my_cos(748)),16);
when x"2ed" => lut_sig <= to_unsigned(integer(my_cos(749)),16);
when x"2ee" => lut_sig <= to_unsigned(integer(my_cos(750)),16);
when x"2ef" => lut_sig <= to_unsigned(integer(my_cos(751)),16);
when x"2f0" => lut_sig <= to_unsigned(integer(my_cos(752)),16);
when x"2f1" => lut_sig <= to_unsigned(integer(my_cos(753)),16);
when x"2f2" => lut_sig <= to_unsigned(integer(my_cos(754)),16);
when x"2f3" => lut_sig <= to_unsigned(integer(my_cos(755)),16);
when x"2f4" => lut_sig <= to_unsigned(integer(my_cos(756)),16);
when x"2f5" => lut_sig <= to_unsigned(integer(my_cos(757)),16);
when x"2f6" => lut_sig <= to_unsigned(integer(my_cos(758)),16);
when x"2f7" => lut_sig <= to_unsigned(integer(my_cos(759)),16);
when x"2f8" => lut_sig <= to_unsigned(integer(my_cos(760)),16);
when x"2f9" => lut_sig <= to_unsigned(integer(my_cos(761)),16);
when x"2fa" => lut_sig <= to_unsigned(integer(my_cos(762)),16);
when x"2fb" => lut_sig <= to_unsigned(integer(my_cos(763)),16);
when x"2fc" => lut_sig <= to_unsigned(integer(my_cos(764)),16);
when x"2fd" => lut_sig <= to_unsigned(integer(my_cos(765)),16);
when x"2fe" => lut_sig <= to_unsigned(integer(my_cos(766)),16);
when x"2ff" => lut_sig <= to_unsigned(integer(my_cos(767)),16);
when x"300" => lut_sig <= to_unsigned(integer(my_cos(768)),16);
when x"301" => lut_sig <= to_unsigned(integer(my_cos(769)),16);
when x"302" => lut_sig <= to_unsigned(integer(my_cos(770)),16);
when x"303" => lut_sig <= to_unsigned(integer(my_cos(771)),16);
when x"304" => lut_sig <= to_unsigned(integer(my_cos(772)),16);
when x"305" => lut_sig <= to_unsigned(integer(my_cos(773)),16);
when x"306" => lut_sig <= to_unsigned(integer(my_cos(774)),16);
when x"307" => lut_sig <= to_unsigned(integer(my_cos(775)),16);
when x"308" => lut_sig <= to_unsigned(integer(my_cos(776)),16);
when x"309" => lut_sig <= to_unsigned(integer(my_cos(777)),16);
when x"30a" => lut_sig <= to_unsigned(integer(my_cos(778)),16);
when x"30b" => lut_sig <= to_unsigned(integer(my_cos(779)),16);
when x"30c" => lut_sig <= to_unsigned(integer(my_cos(780)),16);
when x"30d" => lut_sig <= to_unsigned(integer(my_cos(781)),16);
when x"30e" => lut_sig <= to_unsigned(integer(my_cos(782)),16);
when x"30f" => lut_sig <= to_unsigned(integer(my_cos(783)),16);
when x"310" => lut_sig <= to_unsigned(integer(my_cos(784)),16);
when x"311" => lut_sig <= to_unsigned(integer(my_cos(785)),16);
when x"312" => lut_sig <= to_unsigned(integer(my_cos(786)),16);
when x"313" => lut_sig <= to_unsigned(integer(my_cos(787)),16);
when x"314" => lut_sig <= to_unsigned(integer(my_cos(788)),16);
when x"315" => lut_sig <= to_unsigned(integer(my_cos(789)),16);
when x"316" => lut_sig <= to_unsigned(integer(my_cos(790)),16);
when x"317" => lut_sig <= to_unsigned(integer(my_cos(791)),16);
when x"318" => lut_sig <= to_unsigned(integer(my_cos(792)),16);
when x"319" => lut_sig <= to_unsigned(integer(my_cos(793)),16);
when x"31a" => lut_sig <= to_unsigned(integer(my_cos(794)),16);
when x"31b" => lut_sig <= to_unsigned(integer(my_cos(795)),16);
when x"31c" => lut_sig <= to_unsigned(integer(my_cos(796)),16);
when x"31d" => lut_sig <= to_unsigned(integer(my_cos(797)),16);
when x"31e" => lut_sig <= to_unsigned(integer(my_cos(798)),16);
when x"31f" => lut_sig <= to_unsigned(integer(my_cos(799)),16);
when x"320" => lut_sig <= to_unsigned(integer(my_cos(800)),16);
when x"321" => lut_sig <= to_unsigned(integer(my_cos(801)),16);
when x"322" => lut_sig <= to_unsigned(integer(my_cos(802)),16);
when x"323" => lut_sig <= to_unsigned(integer(my_cos(803)),16);
when x"324" => lut_sig <= to_unsigned(integer(my_cos(804)),16);
when x"325" => lut_sig <= to_unsigned(integer(my_cos(805)),16);
when x"326" => lut_sig <= to_unsigned(integer(my_cos(806)),16);
when x"327" => lut_sig <= to_unsigned(integer(my_cos(807)),16);
when x"328" => lut_sig <= to_unsigned(integer(my_cos(808)),16);
when x"329" => lut_sig <= to_unsigned(integer(my_cos(809)),16);
when x"32a" => lut_sig <= to_unsigned(integer(my_cos(810)),16);
when x"32b" => lut_sig <= to_unsigned(integer(my_cos(811)),16);
when x"32c" => lut_sig <= to_unsigned(integer(my_cos(812)),16);
when x"32d" => lut_sig <= to_unsigned(integer(my_cos(813)),16);
when x"32e" => lut_sig <= to_unsigned(integer(my_cos(814)),16);
when x"32f" => lut_sig <= to_unsigned(integer(my_cos(815)),16);
when x"330" => lut_sig <= to_unsigned(integer(my_cos(816)),16);
when x"331" => lut_sig <= to_unsigned(integer(my_cos(817)),16);
when x"332" => lut_sig <= to_unsigned(integer(my_cos(818)),16);
when x"333" => lut_sig <= to_unsigned(integer(my_cos(819)),16);
when x"334" => lut_sig <= to_unsigned(integer(my_cos(820)),16);
when x"335" => lut_sig <= to_unsigned(integer(my_cos(821)),16);
when x"336" => lut_sig <= to_unsigned(integer(my_cos(822)),16);
when x"337" => lut_sig <= to_unsigned(integer(my_cos(823)),16);
when x"338" => lut_sig <= to_unsigned(integer(my_cos(824)),16);
when x"339" => lut_sig <= to_unsigned(integer(my_cos(825)),16);
when x"33a" => lut_sig <= to_unsigned(integer(my_cos(826)),16);
when x"33b" => lut_sig <= to_unsigned(integer(my_cos(827)),16);
when x"33c" => lut_sig <= to_unsigned(integer(my_cos(828)),16);
when x"33d" => lut_sig <= to_unsigned(integer(my_cos(829)),16);
when x"33e" => lut_sig <= to_unsigned(integer(my_cos(830)),16);
when x"33f" => lut_sig <= to_unsigned(integer(my_cos(831)),16);
when x"340" => lut_sig <= to_unsigned(integer(my_cos(832)),16);
when x"341" => lut_sig <= to_unsigned(integer(my_cos(833)),16);
when x"342" => lut_sig <= to_unsigned(integer(my_cos(834)),16);
when x"343" => lut_sig <= to_unsigned(integer(my_cos(835)),16);
when x"344" => lut_sig <= to_unsigned(integer(my_cos(836)),16);
when x"345" => lut_sig <= to_unsigned(integer(my_cos(837)),16);
when x"346" => lut_sig <= to_unsigned(integer(my_cos(838)),16);
when x"347" => lut_sig <= to_unsigned(integer(my_cos(839)),16);
when x"348" => lut_sig <= to_unsigned(integer(my_cos(840)),16);
when x"349" => lut_sig <= to_unsigned(integer(my_cos(841)),16);
when x"34a" => lut_sig <= to_unsigned(integer(my_cos(842)),16);
when x"34b" => lut_sig <= to_unsigned(integer(my_cos(843)),16);
when x"34c" => lut_sig <= to_unsigned(integer(my_cos(844)),16);
when x"34d" => lut_sig <= to_unsigned(integer(my_cos(845)),16);
when x"34e" => lut_sig <= to_unsigned(integer(my_cos(846)),16);
when x"34f" => lut_sig <= to_unsigned(integer(my_cos(847)),16);
when x"350" => lut_sig <= to_unsigned(integer(my_cos(848)),16);
when x"351" => lut_sig <= to_unsigned(integer(my_cos(849)),16);
when x"352" => lut_sig <= to_unsigned(integer(my_cos(850)),16);
when x"353" => lut_sig <= to_unsigned(integer(my_cos(851)),16);
when x"354" => lut_sig <= to_unsigned(integer(my_cos(852)),16);
when x"355" => lut_sig <= to_unsigned(integer(my_cos(853)),16);
when x"356" => lut_sig <= to_unsigned(integer(my_cos(854)),16);
when x"357" => lut_sig <= to_unsigned(integer(my_cos(855)),16);
when x"358" => lut_sig <= to_unsigned(integer(my_cos(856)),16);
when x"359" => lut_sig <= to_unsigned(integer(my_cos(857)),16);
when x"35a" => lut_sig <= to_unsigned(integer(my_cos(858)),16);
when x"35b" => lut_sig <= to_unsigned(integer(my_cos(859)),16);
when x"35c" => lut_sig <= to_unsigned(integer(my_cos(860)),16);
when x"35d" => lut_sig <= to_unsigned(integer(my_cos(861)),16);
when x"35e" => lut_sig <= to_unsigned(integer(my_cos(862)),16);
when x"35f" => lut_sig <= to_unsigned(integer(my_cos(863)),16);
when x"360" => lut_sig <= to_unsigned(integer(my_cos(864)),16);
when x"361" => lut_sig <= to_unsigned(integer(my_cos(865)),16);
when x"362" => lut_sig <= to_unsigned(integer(my_cos(866)),16);
when x"363" => lut_sig <= to_unsigned(integer(my_cos(867)),16);
when x"364" => lut_sig <= to_unsigned(integer(my_cos(868)),16);
when x"365" => lut_sig <= to_unsigned(integer(my_cos(869)),16);
when x"366" => lut_sig <= to_unsigned(integer(my_cos(870)),16);
when x"367" => lut_sig <= to_unsigned(integer(my_cos(871)),16);
when x"368" => lut_sig <= to_unsigned(integer(my_cos(872)),16);
when x"369" => lut_sig <= to_unsigned(integer(my_cos(873)),16);
when x"36a" => lut_sig <= to_unsigned(integer(my_cos(874)),16);
when x"36b" => lut_sig <= to_unsigned(integer(my_cos(875)),16);
when x"36c" => lut_sig <= to_unsigned(integer(my_cos(876)),16);
when x"36d" => lut_sig <= to_unsigned(integer(my_cos(877)),16);
when x"36e" => lut_sig <= to_unsigned(integer(my_cos(878)),16);
when x"36f" => lut_sig <= to_unsigned(integer(my_cos(879)),16);
when x"370" => lut_sig <= to_unsigned(integer(my_cos(880)),16);
when x"371" => lut_sig <= to_unsigned(integer(my_cos(881)),16);
when x"372" => lut_sig <= to_unsigned(integer(my_cos(882)),16);
when x"373" => lut_sig <= to_unsigned(integer(my_cos(883)),16);
when x"374" => lut_sig <= to_unsigned(integer(my_cos(884)),16);
when x"375" => lut_sig <= to_unsigned(integer(my_cos(885)),16);
when x"376" => lut_sig <= to_unsigned(integer(my_cos(886)),16);
when x"377" => lut_sig <= to_unsigned(integer(my_cos(887)),16);
when x"378" => lut_sig <= to_unsigned(integer(my_cos(888)),16);
when x"379" => lut_sig <= to_unsigned(integer(my_cos(889)),16);
when x"37a" => lut_sig <= to_unsigned(integer(my_cos(890)),16);
when x"37b" => lut_sig <= to_unsigned(integer(my_cos(891)),16);
when x"37c" => lut_sig <= to_unsigned(integer(my_cos(892)),16);
when x"37d" => lut_sig <= to_unsigned(integer(my_cos(893)),16);
when x"37e" => lut_sig <= to_unsigned(integer(my_cos(894)),16);
when x"37f" => lut_sig <= to_unsigned(integer(my_cos(895)),16);
when x"380" => lut_sig <= to_unsigned(integer(my_cos(896)),16);
when x"381" => lut_sig <= to_unsigned(integer(my_cos(897)),16);
when x"382" => lut_sig <= to_unsigned(integer(my_cos(898)),16);
when x"383" => lut_sig <= to_unsigned(integer(my_cos(899)),16);
when x"384" => lut_sig <= to_unsigned(integer(my_cos(900)),16);
when x"385" => lut_sig <= to_unsigned(integer(my_cos(901)),16);
when x"386" => lut_sig <= to_unsigned(integer(my_cos(902)),16);
when x"387" => lut_sig <= to_unsigned(integer(my_cos(903)),16);
when x"388" => lut_sig <= to_unsigned(integer(my_cos(904)),16);
when x"389" => lut_sig <= to_unsigned(integer(my_cos(905)),16);
when x"38a" => lut_sig <= to_unsigned(integer(my_cos(906)),16);
when x"38b" => lut_sig <= to_unsigned(integer(my_cos(907)),16);
when x"38c" => lut_sig <= to_unsigned(integer(my_cos(908)),16);
when x"38d" => lut_sig <= to_unsigned(integer(my_cos(909)),16);
when x"38e" => lut_sig <= to_unsigned(integer(my_cos(910)),16);
when x"38f" => lut_sig <= to_unsigned(integer(my_cos(911)),16);
when x"390" => lut_sig <= to_unsigned(integer(my_cos(912)),16);
when x"391" => lut_sig <= to_unsigned(integer(my_cos(913)),16);
when x"392" => lut_sig <= to_unsigned(integer(my_cos(914)),16);
when x"393" => lut_sig <= to_unsigned(integer(my_cos(915)),16);
when x"394" => lut_sig <= to_unsigned(integer(my_cos(916)),16);
when x"395" => lut_sig <= to_unsigned(integer(my_cos(917)),16);
when x"396" => lut_sig <= to_unsigned(integer(my_cos(918)),16);
when x"397" => lut_sig <= to_unsigned(integer(my_cos(919)),16);
when x"398" => lut_sig <= to_unsigned(integer(my_cos(920)),16);
when x"399" => lut_sig <= to_unsigned(integer(my_cos(921)),16);
when x"39a" => lut_sig <= to_unsigned(integer(my_cos(922)),16);
when x"39b" => lut_sig <= to_unsigned(integer(my_cos(923)),16);
when x"39c" => lut_sig <= to_unsigned(integer(my_cos(924)),16);
when x"39d" => lut_sig <= to_unsigned(integer(my_cos(925)),16);
when x"39e" => lut_sig <= to_unsigned(integer(my_cos(926)),16);
when x"39f" => lut_sig <= to_unsigned(integer(my_cos(927)),16);
when x"3a0" => lut_sig <= to_unsigned(integer(my_cos(928)),16);
when x"3a1" => lut_sig <= to_unsigned(integer(my_cos(929)),16);
when x"3a2" => lut_sig <= to_unsigned(integer(my_cos(930)),16);
when x"3a3" => lut_sig <= to_unsigned(integer(my_cos(931)),16);
when x"3a4" => lut_sig <= to_unsigned(integer(my_cos(932)),16);
when x"3a5" => lut_sig <= to_unsigned(integer(my_cos(933)),16);
when x"3a6" => lut_sig <= to_unsigned(integer(my_cos(934)),16);
when x"3a7" => lut_sig <= to_unsigned(integer(my_cos(935)),16);
when x"3a8" => lut_sig <= to_unsigned(integer(my_cos(936)),16);
when x"3a9" => lut_sig <= to_unsigned(integer(my_cos(937)),16);
when x"3aa" => lut_sig <= to_unsigned(integer(my_cos(938)),16);
when x"3ab" => lut_sig <= to_unsigned(integer(my_cos(939)),16);
when x"3ac" => lut_sig <= to_unsigned(integer(my_cos(940)),16);
when x"3ad" => lut_sig <= to_unsigned(integer(my_cos(941)),16);
when x"3ae" => lut_sig <= to_unsigned(integer(my_cos(942)),16);
when x"3af" => lut_sig <= to_unsigned(integer(my_cos(943)),16);
when x"3b0" => lut_sig <= to_unsigned(integer(my_cos(944)),16);
when x"3b1" => lut_sig <= to_unsigned(integer(my_cos(945)),16);
when x"3b2" => lut_sig <= to_unsigned(integer(my_cos(946)),16);
when x"3b3" => lut_sig <= to_unsigned(integer(my_cos(947)),16);
when x"3b4" => lut_sig <= to_unsigned(integer(my_cos(948)),16);
when x"3b5" => lut_sig <= to_unsigned(integer(my_cos(949)),16);
when x"3b6" => lut_sig <= to_unsigned(integer(my_cos(950)),16);
when x"3b7" => lut_sig <= to_unsigned(integer(my_cos(951)),16);
when x"3b8" => lut_sig <= to_unsigned(integer(my_cos(952)),16);
when x"3b9" => lut_sig <= to_unsigned(integer(my_cos(953)),16);
when x"3ba" => lut_sig <= to_unsigned(integer(my_cos(954)),16);
when x"3bb" => lut_sig <= to_unsigned(integer(my_cos(955)),16);
when x"3bc" => lut_sig <= to_unsigned(integer(my_cos(956)),16);
when x"3bd" => lut_sig <= to_unsigned(integer(my_cos(957)),16);
when x"3be" => lut_sig <= to_unsigned(integer(my_cos(958)),16);
when x"3bf" => lut_sig <= to_unsigned(integer(my_cos(959)),16);
when x"3c0" => lut_sig <= to_unsigned(integer(my_cos(960)),16);
when x"3c1" => lut_sig <= to_unsigned(integer(my_cos(961)),16);
when x"3c2" => lut_sig <= to_unsigned(integer(my_cos(962)),16);
when x"3c3" => lut_sig <= to_unsigned(integer(my_cos(963)),16);
when x"3c4" => lut_sig <= to_unsigned(integer(my_cos(964)),16);
when x"3c5" => lut_sig <= to_unsigned(integer(my_cos(965)),16);
when x"3c6" => lut_sig <= to_unsigned(integer(my_cos(966)),16);
when x"3c7" => lut_sig <= to_unsigned(integer(my_cos(967)),16);
when x"3c8" => lut_sig <= to_unsigned(integer(my_cos(968)),16);
when x"3c9" => lut_sig <= to_unsigned(integer(my_cos(969)),16);
when x"3ca" => lut_sig <= to_unsigned(integer(my_cos(970)),16);
when x"3cb" => lut_sig <= to_unsigned(integer(my_cos(971)),16);
when x"3cc" => lut_sig <= to_unsigned(integer(my_cos(972)),16);
when x"3cd" => lut_sig <= to_unsigned(integer(my_cos(973)),16);
when x"3ce" => lut_sig <= to_unsigned(integer(my_cos(974)),16);
when x"3cf" => lut_sig <= to_unsigned(integer(my_cos(975)),16);
when x"3d0" => lut_sig <= to_unsigned(integer(my_cos(976)),16);
when x"3d1" => lut_sig <= to_unsigned(integer(my_cos(977)),16);
when x"3d2" => lut_sig <= to_unsigned(integer(my_cos(978)),16);
when x"3d3" => lut_sig <= to_unsigned(integer(my_cos(979)),16);
when x"3d4" => lut_sig <= to_unsigned(integer(my_cos(980)),16);
when x"3d5" => lut_sig <= to_unsigned(integer(my_cos(981)),16);
when x"3d6" => lut_sig <= to_unsigned(integer(my_cos(982)),16);
when x"3d7" => lut_sig <= to_unsigned(integer(my_cos(983)),16);
when x"3d8" => lut_sig <= to_unsigned(integer(my_cos(984)),16);
when x"3d9" => lut_sig <= to_unsigned(integer(my_cos(985)),16);
when x"3da" => lut_sig <= to_unsigned(integer(my_cos(986)),16);
when x"3db" => lut_sig <= to_unsigned(integer(my_cos(987)),16);
when x"3dc" => lut_sig <= to_unsigned(integer(my_cos(988)),16);
when x"3dd" => lut_sig <= to_unsigned(integer(my_cos(989)),16);
when x"3de" => lut_sig <= to_unsigned(integer(my_cos(990)),16);
when x"3df" => lut_sig <= to_unsigned(integer(my_cos(991)),16);
when x"3e0" => lut_sig <= to_unsigned(integer(my_cos(992)),16);
when x"3e1" => lut_sig <= to_unsigned(integer(my_cos(993)),16);
when x"3e2" => lut_sig <= to_unsigned(integer(my_cos(994)),16);
when x"3e3" => lut_sig <= to_unsigned(integer(my_cos(995)),16);
when x"3e4" => lut_sig <= to_unsigned(integer(my_cos(996)),16);
when x"3e5" => lut_sig <= to_unsigned(integer(my_cos(997)),16);
when x"3e6" => lut_sig <= to_unsigned(integer(my_cos(998)),16);
when x"3e7" => lut_sig <= to_unsigned(integer(my_cos(999)),16);
when x"3e8" => lut_sig <= to_unsigned(integer(my_cos(1000)),16);
when x"3e9" => lut_sig <= to_unsigned(integer(my_cos(1001)),16);
when x"3ea" => lut_sig <= to_unsigned(integer(my_cos(1002)),16);
when x"3eb" => lut_sig <= to_unsigned(integer(my_cos(1003)),16);
when x"3ec" => lut_sig <= to_unsigned(integer(my_cos(1004)),16);
when x"3ed" => lut_sig <= to_unsigned(integer(my_cos(1005)),16);
when x"3ee" => lut_sig <= to_unsigned(integer(my_cos(1006)),16);
when x"3ef" => lut_sig <= to_unsigned(integer(my_cos(1007)),16);
when x"3f0" => lut_sig <= to_unsigned(integer(my_cos(1008)),16);
when x"3f1" => lut_sig <= to_unsigned(integer(my_cos(1009)),16);
when x"3f2" => lut_sig <= to_unsigned(integer(my_cos(1010)),16);
when x"3f3" => lut_sig <= to_unsigned(integer(my_cos(1011)),16);
when x"3f4" => lut_sig <= to_unsigned(integer(my_cos(1012)),16);
when x"3f5" => lut_sig <= to_unsigned(integer(my_cos(1013)),16);
when x"3f6" => lut_sig <= to_unsigned(integer(my_cos(1014)),16);
when x"3f7" => lut_sig <= to_unsigned(integer(my_cos(1015)),16);
when x"3f8" => lut_sig <= to_unsigned(integer(my_cos(1016)),16);
when x"3f9" => lut_sig <= to_unsigned(integer(my_cos(1017)),16);
when x"3fa" => lut_sig <= to_unsigned(integer(my_cos(1018)),16);
when x"3fb" => lut_sig <= to_unsigned(integer(my_cos(1019)),16);
when x"3fc" => lut_sig <= to_unsigned(integer(my_cos(1020)),16);
when x"3fd" => lut_sig <= to_unsigned(integer(my_cos(1021)),16);
when x"3fe" => lut_sig <= to_unsigned(integer(my_cos(1022)),16);
when x"3ff" => lut_sig <= to_unsigned(integer(my_cos(1023)),16);
when x"400" => lut_sig <= to_unsigned(integer(my_cos(1024)),16);
when x"401" => lut_sig <= to_unsigned(integer(my_cos(1025)),16);
when x"402" => lut_sig <= to_unsigned(integer(my_cos(1026)),16);
when x"403" => lut_sig <= to_unsigned(integer(my_cos(1027)),16);
when x"404" => lut_sig <= to_unsigned(integer(my_cos(1028)),16);
when x"405" => lut_sig <= to_unsigned(integer(my_cos(1029)),16);
when x"406" => lut_sig <= to_unsigned(integer(my_cos(1030)),16);
when x"407" => lut_sig <= to_unsigned(integer(my_cos(1031)),16);
when x"408" => lut_sig <= to_unsigned(integer(my_cos(1032)),16);
when x"409" => lut_sig <= to_unsigned(integer(my_cos(1033)),16);
when x"40a" => lut_sig <= to_unsigned(integer(my_cos(1034)),16);
when x"40b" => lut_sig <= to_unsigned(integer(my_cos(1035)),16);
when x"40c" => lut_sig <= to_unsigned(integer(my_cos(1036)),16);
when x"40d" => lut_sig <= to_unsigned(integer(my_cos(1037)),16);
when x"40e" => lut_sig <= to_unsigned(integer(my_cos(1038)),16);
when x"40f" => lut_sig <= to_unsigned(integer(my_cos(1039)),16);
when x"410" => lut_sig <= to_unsigned(integer(my_cos(1040)),16);
when x"411" => lut_sig <= to_unsigned(integer(my_cos(1041)),16);
when x"412" => lut_sig <= to_unsigned(integer(my_cos(1042)),16);
when x"413" => lut_sig <= to_unsigned(integer(my_cos(1043)),16);
when x"414" => lut_sig <= to_unsigned(integer(my_cos(1044)),16);
when x"415" => lut_sig <= to_unsigned(integer(my_cos(1045)),16);
when x"416" => lut_sig <= to_unsigned(integer(my_cos(1046)),16);
when x"417" => lut_sig <= to_unsigned(integer(my_cos(1047)),16);
when x"418" => lut_sig <= to_unsigned(integer(my_cos(1048)),16);
when x"419" => lut_sig <= to_unsigned(integer(my_cos(1049)),16);
when x"41a" => lut_sig <= to_unsigned(integer(my_cos(1050)),16);
when x"41b" => lut_sig <= to_unsigned(integer(my_cos(1051)),16);
when x"41c" => lut_sig <= to_unsigned(integer(my_cos(1052)),16);
when x"41d" => lut_sig <= to_unsigned(integer(my_cos(1053)),16);
when x"41e" => lut_sig <= to_unsigned(integer(my_cos(1054)),16);
when x"41f" => lut_sig <= to_unsigned(integer(my_cos(1055)),16);
when x"420" => lut_sig <= to_unsigned(integer(my_cos(1056)),16);
when x"421" => lut_sig <= to_unsigned(integer(my_cos(1057)),16);
when x"422" => lut_sig <= to_unsigned(integer(my_cos(1058)),16);
when x"423" => lut_sig <= to_unsigned(integer(my_cos(1059)),16);
when x"424" => lut_sig <= to_unsigned(integer(my_cos(1060)),16);
when x"425" => lut_sig <= to_unsigned(integer(my_cos(1061)),16);
when x"426" => lut_sig <= to_unsigned(integer(my_cos(1062)),16);
when x"427" => lut_sig <= to_unsigned(integer(my_cos(1063)),16);
when x"428" => lut_sig <= to_unsigned(integer(my_cos(1064)),16);
when x"429" => lut_sig <= to_unsigned(integer(my_cos(1065)),16);
when x"42a" => lut_sig <= to_unsigned(integer(my_cos(1066)),16);
when x"42b" => lut_sig <= to_unsigned(integer(my_cos(1067)),16);
when x"42c" => lut_sig <= to_unsigned(integer(my_cos(1068)),16);
when x"42d" => lut_sig <= to_unsigned(integer(my_cos(1069)),16);
when x"42e" => lut_sig <= to_unsigned(integer(my_cos(1070)),16);
when x"42f" => lut_sig <= to_unsigned(integer(my_cos(1071)),16);
when x"430" => lut_sig <= to_unsigned(integer(my_cos(1072)),16);
when x"431" => lut_sig <= to_unsigned(integer(my_cos(1073)),16);
when x"432" => lut_sig <= to_unsigned(integer(my_cos(1074)),16);
when x"433" => lut_sig <= to_unsigned(integer(my_cos(1075)),16);
when x"434" => lut_sig <= to_unsigned(integer(my_cos(1076)),16);
when x"435" => lut_sig <= to_unsigned(integer(my_cos(1077)),16);
when x"436" => lut_sig <= to_unsigned(integer(my_cos(1078)),16);
when x"437" => lut_sig <= to_unsigned(integer(my_cos(1079)),16);
when x"438" => lut_sig <= to_unsigned(integer(my_cos(1080)),16);
when x"439" => lut_sig <= to_unsigned(integer(my_cos(1081)),16);
when x"43a" => lut_sig <= to_unsigned(integer(my_cos(1082)),16);
when x"43b" => lut_sig <= to_unsigned(integer(my_cos(1083)),16);
when x"43c" => lut_sig <= to_unsigned(integer(my_cos(1084)),16);
when x"43d" => lut_sig <= to_unsigned(integer(my_cos(1085)),16);
when x"43e" => lut_sig <= to_unsigned(integer(my_cos(1086)),16);
when x"43f" => lut_sig <= to_unsigned(integer(my_cos(1087)),16);
when x"440" => lut_sig <= to_unsigned(integer(my_cos(1088)),16);
when x"441" => lut_sig <= to_unsigned(integer(my_cos(1089)),16);
when x"442" => lut_sig <= to_unsigned(integer(my_cos(1090)),16);
when x"443" => lut_sig <= to_unsigned(integer(my_cos(1091)),16);
when x"444" => lut_sig <= to_unsigned(integer(my_cos(1092)),16);
when x"445" => lut_sig <= to_unsigned(integer(my_cos(1093)),16);
when x"446" => lut_sig <= to_unsigned(integer(my_cos(1094)),16);
when x"447" => lut_sig <= to_unsigned(integer(my_cos(1095)),16);
when x"448" => lut_sig <= to_unsigned(integer(my_cos(1096)),16);
when x"449" => lut_sig <= to_unsigned(integer(my_cos(1097)),16);
when x"44a" => lut_sig <= to_unsigned(integer(my_cos(1098)),16);
when x"44b" => lut_sig <= to_unsigned(integer(my_cos(1099)),16);
when x"44c" => lut_sig <= to_unsigned(integer(my_cos(1100)),16);
when x"44d" => lut_sig <= to_unsigned(integer(my_cos(1101)),16);
when x"44e" => lut_sig <= to_unsigned(integer(my_cos(1102)),16);
when x"44f" => lut_sig <= to_unsigned(integer(my_cos(1103)),16);
when x"450" => lut_sig <= to_unsigned(integer(my_cos(1104)),16);
when x"451" => lut_sig <= to_unsigned(integer(my_cos(1105)),16);
when x"452" => lut_sig <= to_unsigned(integer(my_cos(1106)),16);
when x"453" => lut_sig <= to_unsigned(integer(my_cos(1107)),16);
when x"454" => lut_sig <= to_unsigned(integer(my_cos(1108)),16);
when x"455" => lut_sig <= to_unsigned(integer(my_cos(1109)),16);
when x"456" => lut_sig <= to_unsigned(integer(my_cos(1110)),16);
when x"457" => lut_sig <= to_unsigned(integer(my_cos(1111)),16);
when x"458" => lut_sig <= to_unsigned(integer(my_cos(1112)),16);
when x"459" => lut_sig <= to_unsigned(integer(my_cos(1113)),16);
when x"45a" => lut_sig <= to_unsigned(integer(my_cos(1114)),16);
when x"45b" => lut_sig <= to_unsigned(integer(my_cos(1115)),16);
when x"45c" => lut_sig <= to_unsigned(integer(my_cos(1116)),16);
when x"45d" => lut_sig <= to_unsigned(integer(my_cos(1117)),16);
when x"45e" => lut_sig <= to_unsigned(integer(my_cos(1118)),16);
when x"45f" => lut_sig <= to_unsigned(integer(my_cos(1119)),16);
when x"460" => lut_sig <= to_unsigned(integer(my_cos(1120)),16);
when x"461" => lut_sig <= to_unsigned(integer(my_cos(1121)),16);
when x"462" => lut_sig <= to_unsigned(integer(my_cos(1122)),16);
when x"463" => lut_sig <= to_unsigned(integer(my_cos(1123)),16);
when x"464" => lut_sig <= to_unsigned(integer(my_cos(1124)),16);
when x"465" => lut_sig <= to_unsigned(integer(my_cos(1125)),16);
when x"466" => lut_sig <= to_unsigned(integer(my_cos(1126)),16);
when x"467" => lut_sig <= to_unsigned(integer(my_cos(1127)),16);
when x"468" => lut_sig <= to_unsigned(integer(my_cos(1128)),16);
when x"469" => lut_sig <= to_unsigned(integer(my_cos(1129)),16);
when x"46a" => lut_sig <= to_unsigned(integer(my_cos(1130)),16);
when x"46b" => lut_sig <= to_unsigned(integer(my_cos(1131)),16);
when x"46c" => lut_sig <= to_unsigned(integer(my_cos(1132)),16);
when x"46d" => lut_sig <= to_unsigned(integer(my_cos(1133)),16);
when x"46e" => lut_sig <= to_unsigned(integer(my_cos(1134)),16);
when x"46f" => lut_sig <= to_unsigned(integer(my_cos(1135)),16);
when x"470" => lut_sig <= to_unsigned(integer(my_cos(1136)),16);
when x"471" => lut_sig <= to_unsigned(integer(my_cos(1137)),16);
when x"472" => lut_sig <= to_unsigned(integer(my_cos(1138)),16);
when x"473" => lut_sig <= to_unsigned(integer(my_cos(1139)),16);
when x"474" => lut_sig <= to_unsigned(integer(my_cos(1140)),16);
when x"475" => lut_sig <= to_unsigned(integer(my_cos(1141)),16);
when x"476" => lut_sig <= to_unsigned(integer(my_cos(1142)),16);
when x"477" => lut_sig <= to_unsigned(integer(my_cos(1143)),16);
when x"478" => lut_sig <= to_unsigned(integer(my_cos(1144)),16);
when x"479" => lut_sig <= to_unsigned(integer(my_cos(1145)),16);
when x"47a" => lut_sig <= to_unsigned(integer(my_cos(1146)),16);
when x"47b" => lut_sig <= to_unsigned(integer(my_cos(1147)),16);
when x"47c" => lut_sig <= to_unsigned(integer(my_cos(1148)),16);
when x"47d" => lut_sig <= to_unsigned(integer(my_cos(1149)),16);
when x"47e" => lut_sig <= to_unsigned(integer(my_cos(1150)),16);
when x"47f" => lut_sig <= to_unsigned(integer(my_cos(1151)),16);
when x"480" => lut_sig <= to_unsigned(integer(my_cos(1152)),16);
when x"481" => lut_sig <= to_unsigned(integer(my_cos(1153)),16);
when x"482" => lut_sig <= to_unsigned(integer(my_cos(1154)),16);
when x"483" => lut_sig <= to_unsigned(integer(my_cos(1155)),16);
when x"484" => lut_sig <= to_unsigned(integer(my_cos(1156)),16);
when x"485" => lut_sig <= to_unsigned(integer(my_cos(1157)),16);
when x"486" => lut_sig <= to_unsigned(integer(my_cos(1158)),16);
when x"487" => lut_sig <= to_unsigned(integer(my_cos(1159)),16);
when x"488" => lut_sig <= to_unsigned(integer(my_cos(1160)),16);
when x"489" => lut_sig <= to_unsigned(integer(my_cos(1161)),16);
when x"48a" => lut_sig <= to_unsigned(integer(my_cos(1162)),16);
when x"48b" => lut_sig <= to_unsigned(integer(my_cos(1163)),16);
when x"48c" => lut_sig <= to_unsigned(integer(my_cos(1164)),16);
when x"48d" => lut_sig <= to_unsigned(integer(my_cos(1165)),16);
when x"48e" => lut_sig <= to_unsigned(integer(my_cos(1166)),16);
when x"48f" => lut_sig <= to_unsigned(integer(my_cos(1167)),16);
when x"490" => lut_sig <= to_unsigned(integer(my_cos(1168)),16);
when x"491" => lut_sig <= to_unsigned(integer(my_cos(1169)),16);
when x"492" => lut_sig <= to_unsigned(integer(my_cos(1170)),16);
when x"493" => lut_sig <= to_unsigned(integer(my_cos(1171)),16);
when x"494" => lut_sig <= to_unsigned(integer(my_cos(1172)),16);
when x"495" => lut_sig <= to_unsigned(integer(my_cos(1173)),16);
when x"496" => lut_sig <= to_unsigned(integer(my_cos(1174)),16);
when x"497" => lut_sig <= to_unsigned(integer(my_cos(1175)),16);
when x"498" => lut_sig <= to_unsigned(integer(my_cos(1176)),16);
when x"499" => lut_sig <= to_unsigned(integer(my_cos(1177)),16);
when x"49a" => lut_sig <= to_unsigned(integer(my_cos(1178)),16);
when x"49b" => lut_sig <= to_unsigned(integer(my_cos(1179)),16);
when x"49c" => lut_sig <= to_unsigned(integer(my_cos(1180)),16);
when x"49d" => lut_sig <= to_unsigned(integer(my_cos(1181)),16);
when x"49e" => lut_sig <= to_unsigned(integer(my_cos(1182)),16);
when x"49f" => lut_sig <= to_unsigned(integer(my_cos(1183)),16);
when x"4a0" => lut_sig <= to_unsigned(integer(my_cos(1184)),16);
when x"4a1" => lut_sig <= to_unsigned(integer(my_cos(1185)),16);
when x"4a2" => lut_sig <= to_unsigned(integer(my_cos(1186)),16);
when x"4a3" => lut_sig <= to_unsigned(integer(my_cos(1187)),16);
when x"4a4" => lut_sig <= to_unsigned(integer(my_cos(1188)),16);
when x"4a5" => lut_sig <= to_unsigned(integer(my_cos(1189)),16);
when x"4a6" => lut_sig <= to_unsigned(integer(my_cos(1190)),16);
when x"4a7" => lut_sig <= to_unsigned(integer(my_cos(1191)),16);
when x"4a8" => lut_sig <= to_unsigned(integer(my_cos(1192)),16);
when x"4a9" => lut_sig <= to_unsigned(integer(my_cos(1193)),16);
when x"4aa" => lut_sig <= to_unsigned(integer(my_cos(1194)),16);
when x"4ab" => lut_sig <= to_unsigned(integer(my_cos(1195)),16);
when x"4ac" => lut_sig <= to_unsigned(integer(my_cos(1196)),16);
when x"4ad" => lut_sig <= to_unsigned(integer(my_cos(1197)),16);
when x"4ae" => lut_sig <= to_unsigned(integer(my_cos(1198)),16);
when x"4af" => lut_sig <= to_unsigned(integer(my_cos(1199)),16);
when x"4b0" => lut_sig <= to_unsigned(integer(my_cos(1200)),16);
when x"4b1" => lut_sig <= to_unsigned(integer(my_cos(1201)),16);
when x"4b2" => lut_sig <= to_unsigned(integer(my_cos(1202)),16);
when x"4b3" => lut_sig <= to_unsigned(integer(my_cos(1203)),16);
when x"4b4" => lut_sig <= to_unsigned(integer(my_cos(1204)),16);
when x"4b5" => lut_sig <= to_unsigned(integer(my_cos(1205)),16);
when x"4b6" => lut_sig <= to_unsigned(integer(my_cos(1206)),16);
when x"4b7" => lut_sig <= to_unsigned(integer(my_cos(1207)),16);
when x"4b8" => lut_sig <= to_unsigned(integer(my_cos(1208)),16);
when x"4b9" => lut_sig <= to_unsigned(integer(my_cos(1209)),16);
when x"4ba" => lut_sig <= to_unsigned(integer(my_cos(1210)),16);
when x"4bb" => lut_sig <= to_unsigned(integer(my_cos(1211)),16);
when x"4bc" => lut_sig <= to_unsigned(integer(my_cos(1212)),16);
when x"4bd" => lut_sig <= to_unsigned(integer(my_cos(1213)),16);
when x"4be" => lut_sig <= to_unsigned(integer(my_cos(1214)),16);
when x"4bf" => lut_sig <= to_unsigned(integer(my_cos(1215)),16);
when x"4c0" => lut_sig <= to_unsigned(integer(my_cos(1216)),16);
when x"4c1" => lut_sig <= to_unsigned(integer(my_cos(1217)),16);
when x"4c2" => lut_sig <= to_unsigned(integer(my_cos(1218)),16);
when x"4c3" => lut_sig <= to_unsigned(integer(my_cos(1219)),16);
when x"4c4" => lut_sig <= to_unsigned(integer(my_cos(1220)),16);
when x"4c5" => lut_sig <= to_unsigned(integer(my_cos(1221)),16);
when x"4c6" => lut_sig <= to_unsigned(integer(my_cos(1222)),16);
when x"4c7" => lut_sig <= to_unsigned(integer(my_cos(1223)),16);
when x"4c8" => lut_sig <= to_unsigned(integer(my_cos(1224)),16);
when x"4c9" => lut_sig <= to_unsigned(integer(my_cos(1225)),16);
when x"4ca" => lut_sig <= to_unsigned(integer(my_cos(1226)),16);
when x"4cb" => lut_sig <= to_unsigned(integer(my_cos(1227)),16);
when x"4cc" => lut_sig <= to_unsigned(integer(my_cos(1228)),16);
when x"4cd" => lut_sig <= to_unsigned(integer(my_cos(1229)),16);
when x"4ce" => lut_sig <= to_unsigned(integer(my_cos(1230)),16);
when x"4cf" => lut_sig <= to_unsigned(integer(my_cos(1231)),16);
when x"4d0" => lut_sig <= to_unsigned(integer(my_cos(1232)),16);
when x"4d1" => lut_sig <= to_unsigned(integer(my_cos(1233)),16);
when x"4d2" => lut_sig <= to_unsigned(integer(my_cos(1234)),16);
when x"4d3" => lut_sig <= to_unsigned(integer(my_cos(1235)),16);
when x"4d4" => lut_sig <= to_unsigned(integer(my_cos(1236)),16);
when x"4d5" => lut_sig <= to_unsigned(integer(my_cos(1237)),16);
when x"4d6" => lut_sig <= to_unsigned(integer(my_cos(1238)),16);
when x"4d7" => lut_sig <= to_unsigned(integer(my_cos(1239)),16);
when x"4d8" => lut_sig <= to_unsigned(integer(my_cos(1240)),16);
when x"4d9" => lut_sig <= to_unsigned(integer(my_cos(1241)),16);
when x"4da" => lut_sig <= to_unsigned(integer(my_cos(1242)),16);
when x"4db" => lut_sig <= to_unsigned(integer(my_cos(1243)),16);
when x"4dc" => lut_sig <= to_unsigned(integer(my_cos(1244)),16);
when x"4dd" => lut_sig <= to_unsigned(integer(my_cos(1245)),16);
when x"4de" => lut_sig <= to_unsigned(integer(my_cos(1246)),16);
when x"4df" => lut_sig <= to_unsigned(integer(my_cos(1247)),16);
when x"4e0" => lut_sig <= to_unsigned(integer(my_cos(1248)),16);
when x"4e1" => lut_sig <= to_unsigned(integer(my_cos(1249)),16);
when x"4e2" => lut_sig <= to_unsigned(integer(my_cos(1250)),16);
when x"4e3" => lut_sig <= to_unsigned(integer(my_cos(1251)),16);
when x"4e4" => lut_sig <= to_unsigned(integer(my_cos(1252)),16);
when x"4e5" => lut_sig <= to_unsigned(integer(my_cos(1253)),16);
when x"4e6" => lut_sig <= to_unsigned(integer(my_cos(1254)),16);
when x"4e7" => lut_sig <= to_unsigned(integer(my_cos(1255)),16);
when x"4e8" => lut_sig <= to_unsigned(integer(my_cos(1256)),16);
when x"4e9" => lut_sig <= to_unsigned(integer(my_cos(1257)),16);
when x"4ea" => lut_sig <= to_unsigned(integer(my_cos(1258)),16);
when x"4eb" => lut_sig <= to_unsigned(integer(my_cos(1259)),16);
when x"4ec" => lut_sig <= to_unsigned(integer(my_cos(1260)),16);
when x"4ed" => lut_sig <= to_unsigned(integer(my_cos(1261)),16);
when x"4ee" => lut_sig <= to_unsigned(integer(my_cos(1262)),16);
when x"4ef" => lut_sig <= to_unsigned(integer(my_cos(1263)),16);
when x"4f0" => lut_sig <= to_unsigned(integer(my_cos(1264)),16);
when x"4f1" => lut_sig <= to_unsigned(integer(my_cos(1265)),16);
when x"4f2" => lut_sig <= to_unsigned(integer(my_cos(1266)),16);
when x"4f3" => lut_sig <= to_unsigned(integer(my_cos(1267)),16);
when x"4f4" => lut_sig <= to_unsigned(integer(my_cos(1268)),16);
when x"4f5" => lut_sig <= to_unsigned(integer(my_cos(1269)),16);
when x"4f6" => lut_sig <= to_unsigned(integer(my_cos(1270)),16);
when x"4f7" => lut_sig <= to_unsigned(integer(my_cos(1271)),16);
when x"4f8" => lut_sig <= to_unsigned(integer(my_cos(1272)),16);
when x"4f9" => lut_sig <= to_unsigned(integer(my_cos(1273)),16);
when x"4fa" => lut_sig <= to_unsigned(integer(my_cos(1274)),16);
when x"4fb" => lut_sig <= to_unsigned(integer(my_cos(1275)),16);
when x"4fc" => lut_sig <= to_unsigned(integer(my_cos(1276)),16);
when x"4fd" => lut_sig <= to_unsigned(integer(my_cos(1277)),16);
when x"4fe" => lut_sig <= to_unsigned(integer(my_cos(1278)),16);
when x"4ff" => lut_sig <= to_unsigned(integer(my_cos(1279)),16);
when x"500" => lut_sig <= to_unsigned(integer(my_cos(1280)),16);
when x"501" => lut_sig <= to_unsigned(integer(my_cos(1281)),16);
when x"502" => lut_sig <= to_unsigned(integer(my_cos(1282)),16);
when x"503" => lut_sig <= to_unsigned(integer(my_cos(1283)),16);
when x"504" => lut_sig <= to_unsigned(integer(my_cos(1284)),16);
when x"505" => lut_sig <= to_unsigned(integer(my_cos(1285)),16);
when x"506" => lut_sig <= to_unsigned(integer(my_cos(1286)),16);
when x"507" => lut_sig <= to_unsigned(integer(my_cos(1287)),16);
when x"508" => lut_sig <= to_unsigned(integer(my_cos(1288)),16);
when x"509" => lut_sig <= to_unsigned(integer(my_cos(1289)),16);
when x"50a" => lut_sig <= to_unsigned(integer(my_cos(1290)),16);
when x"50b" => lut_sig <= to_unsigned(integer(my_cos(1291)),16);
when x"50c" => lut_sig <= to_unsigned(integer(my_cos(1292)),16);
when x"50d" => lut_sig <= to_unsigned(integer(my_cos(1293)),16);
when x"50e" => lut_sig <= to_unsigned(integer(my_cos(1294)),16);
when x"50f" => lut_sig <= to_unsigned(integer(my_cos(1295)),16);
when x"510" => lut_sig <= to_unsigned(integer(my_cos(1296)),16);
when x"511" => lut_sig <= to_unsigned(integer(my_cos(1297)),16);
when x"512" => lut_sig <= to_unsigned(integer(my_cos(1298)),16);
when x"513" => lut_sig <= to_unsigned(integer(my_cos(1299)),16);
when x"514" => lut_sig <= to_unsigned(integer(my_cos(1300)),16);
when x"515" => lut_sig <= to_unsigned(integer(my_cos(1301)),16);
when x"516" => lut_sig <= to_unsigned(integer(my_cos(1302)),16);
when x"517" => lut_sig <= to_unsigned(integer(my_cos(1303)),16);
when x"518" => lut_sig <= to_unsigned(integer(my_cos(1304)),16);
when x"519" => lut_sig <= to_unsigned(integer(my_cos(1305)),16);
when x"51a" => lut_sig <= to_unsigned(integer(my_cos(1306)),16);
when x"51b" => lut_sig <= to_unsigned(integer(my_cos(1307)),16);
when x"51c" => lut_sig <= to_unsigned(integer(my_cos(1308)),16);
when x"51d" => lut_sig <= to_unsigned(integer(my_cos(1309)),16);
when x"51e" => lut_sig <= to_unsigned(integer(my_cos(1310)),16);
when x"51f" => lut_sig <= to_unsigned(integer(my_cos(1311)),16);
when x"520" => lut_sig <= to_unsigned(integer(my_cos(1312)),16);
when x"521" => lut_sig <= to_unsigned(integer(my_cos(1313)),16);
when x"522" => lut_sig <= to_unsigned(integer(my_cos(1314)),16);
when x"523" => lut_sig <= to_unsigned(integer(my_cos(1315)),16);
when x"524" => lut_sig <= to_unsigned(integer(my_cos(1316)),16);
when x"525" => lut_sig <= to_unsigned(integer(my_cos(1317)),16);
when x"526" => lut_sig <= to_unsigned(integer(my_cos(1318)),16);
when x"527" => lut_sig <= to_unsigned(integer(my_cos(1319)),16);
when x"528" => lut_sig <= to_unsigned(integer(my_cos(1320)),16);
when x"529" => lut_sig <= to_unsigned(integer(my_cos(1321)),16);
when x"52a" => lut_sig <= to_unsigned(integer(my_cos(1322)),16);
when x"52b" => lut_sig <= to_unsigned(integer(my_cos(1323)),16);
when x"52c" => lut_sig <= to_unsigned(integer(my_cos(1324)),16);
when x"52d" => lut_sig <= to_unsigned(integer(my_cos(1325)),16);
when x"52e" => lut_sig <= to_unsigned(integer(my_cos(1326)),16);
when x"52f" => lut_sig <= to_unsigned(integer(my_cos(1327)),16);
when x"530" => lut_sig <= to_unsigned(integer(my_cos(1328)),16);
when x"531" => lut_sig <= to_unsigned(integer(my_cos(1329)),16);
when x"532" => lut_sig <= to_unsigned(integer(my_cos(1330)),16);
when x"533" => lut_sig <= to_unsigned(integer(my_cos(1331)),16);
when x"534" => lut_sig <= to_unsigned(integer(my_cos(1332)),16);
when x"535" => lut_sig <= to_unsigned(integer(my_cos(1333)),16);
when x"536" => lut_sig <= to_unsigned(integer(my_cos(1334)),16);
when x"537" => lut_sig <= to_unsigned(integer(my_cos(1335)),16);
when x"538" => lut_sig <= to_unsigned(integer(my_cos(1336)),16);
when x"539" => lut_sig <= to_unsigned(integer(my_cos(1337)),16);
when x"53a" => lut_sig <= to_unsigned(integer(my_cos(1338)),16);
when x"53b" => lut_sig <= to_unsigned(integer(my_cos(1339)),16);
when x"53c" => lut_sig <= to_unsigned(integer(my_cos(1340)),16);
when x"53d" => lut_sig <= to_unsigned(integer(my_cos(1341)),16);
when x"53e" => lut_sig <= to_unsigned(integer(my_cos(1342)),16);
when x"53f" => lut_sig <= to_unsigned(integer(my_cos(1343)),16);
when x"540" => lut_sig <= to_unsigned(integer(my_cos(1344)),16);
when x"541" => lut_sig <= to_unsigned(integer(my_cos(1345)),16);
when x"542" => lut_sig <= to_unsigned(integer(my_cos(1346)),16);
when x"543" => lut_sig <= to_unsigned(integer(my_cos(1347)),16);
when x"544" => lut_sig <= to_unsigned(integer(my_cos(1348)),16);
when x"545" => lut_sig <= to_unsigned(integer(my_cos(1349)),16);
when x"546" => lut_sig <= to_unsigned(integer(my_cos(1350)),16);
when x"547" => lut_sig <= to_unsigned(integer(my_cos(1351)),16);
when x"548" => lut_sig <= to_unsigned(integer(my_cos(1352)),16);
when x"549" => lut_sig <= to_unsigned(integer(my_cos(1353)),16);
when x"54a" => lut_sig <= to_unsigned(integer(my_cos(1354)),16);
when x"54b" => lut_sig <= to_unsigned(integer(my_cos(1355)),16);
when x"54c" => lut_sig <= to_unsigned(integer(my_cos(1356)),16);
when x"54d" => lut_sig <= to_unsigned(integer(my_cos(1357)),16);
when x"54e" => lut_sig <= to_unsigned(integer(my_cos(1358)),16);
when x"54f" => lut_sig <= to_unsigned(integer(my_cos(1359)),16);
when x"550" => lut_sig <= to_unsigned(integer(my_cos(1360)),16);
when x"551" => lut_sig <= to_unsigned(integer(my_cos(1361)),16);
when x"552" => lut_sig <= to_unsigned(integer(my_cos(1362)),16);
when x"553" => lut_sig <= to_unsigned(integer(my_cos(1363)),16);
when x"554" => lut_sig <= to_unsigned(integer(my_cos(1364)),16);
when x"555" => lut_sig <= to_unsigned(integer(my_cos(1365)),16);
when x"556" => lut_sig <= to_unsigned(integer(my_cos(1366)),16);
when x"557" => lut_sig <= to_unsigned(integer(my_cos(1367)),16);
when x"558" => lut_sig <= to_unsigned(integer(my_cos(1368)),16);
when x"559" => lut_sig <= to_unsigned(integer(my_cos(1369)),16);
when x"55a" => lut_sig <= to_unsigned(integer(my_cos(1370)),16);
when x"55b" => lut_sig <= to_unsigned(integer(my_cos(1371)),16);
when x"55c" => lut_sig <= to_unsigned(integer(my_cos(1372)),16);
when x"55d" => lut_sig <= to_unsigned(integer(my_cos(1373)),16);
when x"55e" => lut_sig <= to_unsigned(integer(my_cos(1374)),16);
when x"55f" => lut_sig <= to_unsigned(integer(my_cos(1375)),16);
when x"560" => lut_sig <= to_unsigned(integer(my_cos(1376)),16);
when x"561" => lut_sig <= to_unsigned(integer(my_cos(1377)),16);
when x"562" => lut_sig <= to_unsigned(integer(my_cos(1378)),16);
when x"563" => lut_sig <= to_unsigned(integer(my_cos(1379)),16);
when x"564" => lut_sig <= to_unsigned(integer(my_cos(1380)),16);
when x"565" => lut_sig <= to_unsigned(integer(my_cos(1381)),16);
when x"566" => lut_sig <= to_unsigned(integer(my_cos(1382)),16);
when x"567" => lut_sig <= to_unsigned(integer(my_cos(1383)),16);
when x"568" => lut_sig <= to_unsigned(integer(my_cos(1384)),16);
when x"569" => lut_sig <= to_unsigned(integer(my_cos(1385)),16);
when x"56a" => lut_sig <= to_unsigned(integer(my_cos(1386)),16);
when x"56b" => lut_sig <= to_unsigned(integer(my_cos(1387)),16);
when x"56c" => lut_sig <= to_unsigned(integer(my_cos(1388)),16);
when x"56d" => lut_sig <= to_unsigned(integer(my_cos(1389)),16);
when x"56e" => lut_sig <= to_unsigned(integer(my_cos(1390)),16);
when x"56f" => lut_sig <= to_unsigned(integer(my_cos(1391)),16);
when x"570" => lut_sig <= to_unsigned(integer(my_cos(1392)),16);
when x"571" => lut_sig <= to_unsigned(integer(my_cos(1393)),16);
when x"572" => lut_sig <= to_unsigned(integer(my_cos(1394)),16);
when x"573" => lut_sig <= to_unsigned(integer(my_cos(1395)),16);
when x"574" => lut_sig <= to_unsigned(integer(my_cos(1396)),16);
when x"575" => lut_sig <= to_unsigned(integer(my_cos(1397)),16);
when x"576" => lut_sig <= to_unsigned(integer(my_cos(1398)),16);
when x"577" => lut_sig <= to_unsigned(integer(my_cos(1399)),16);
when x"578" => lut_sig <= to_unsigned(integer(my_cos(1400)),16);
when x"579" => lut_sig <= to_unsigned(integer(my_cos(1401)),16);
when x"57a" => lut_sig <= to_unsigned(integer(my_cos(1402)),16);
when x"57b" => lut_sig <= to_unsigned(integer(my_cos(1403)),16);
when x"57c" => lut_sig <= to_unsigned(integer(my_cos(1404)),16);
when x"57d" => lut_sig <= to_unsigned(integer(my_cos(1405)),16);
when x"57e" => lut_sig <= to_unsigned(integer(my_cos(1406)),16);
when x"57f" => lut_sig <= to_unsigned(integer(my_cos(1407)),16);
when x"580" => lut_sig <= to_unsigned(integer(my_cos(1408)),16);
when x"581" => lut_sig <= to_unsigned(integer(my_cos(1409)),16);
when x"582" => lut_sig <= to_unsigned(integer(my_cos(1410)),16);
when x"583" => lut_sig <= to_unsigned(integer(my_cos(1411)),16);
when x"584" => lut_sig <= to_unsigned(integer(my_cos(1412)),16);
when x"585" => lut_sig <= to_unsigned(integer(my_cos(1413)),16);
when x"586" => lut_sig <= to_unsigned(integer(my_cos(1414)),16);
when x"587" => lut_sig <= to_unsigned(integer(my_cos(1415)),16);
when x"588" => lut_sig <= to_unsigned(integer(my_cos(1416)),16);
when x"589" => lut_sig <= to_unsigned(integer(my_cos(1417)),16);
when x"58a" => lut_sig <= to_unsigned(integer(my_cos(1418)),16);
when x"58b" => lut_sig <= to_unsigned(integer(my_cos(1419)),16);
when x"58c" => lut_sig <= to_unsigned(integer(my_cos(1420)),16);
when x"58d" => lut_sig <= to_unsigned(integer(my_cos(1421)),16);
when x"58e" => lut_sig <= to_unsigned(integer(my_cos(1422)),16);
when x"58f" => lut_sig <= to_unsigned(integer(my_cos(1423)),16);
when x"590" => lut_sig <= to_unsigned(integer(my_cos(1424)),16);
when x"591" => lut_sig <= to_unsigned(integer(my_cos(1425)),16);
when x"592" => lut_sig <= to_unsigned(integer(my_cos(1426)),16);
when x"593" => lut_sig <= to_unsigned(integer(my_cos(1427)),16);
when x"594" => lut_sig <= to_unsigned(integer(my_cos(1428)),16);
when x"595" => lut_sig <= to_unsigned(integer(my_cos(1429)),16);
when x"596" => lut_sig <= to_unsigned(integer(my_cos(1430)),16);
when x"597" => lut_sig <= to_unsigned(integer(my_cos(1431)),16);
when x"598" => lut_sig <= to_unsigned(integer(my_cos(1432)),16);
when x"599" => lut_sig <= to_unsigned(integer(my_cos(1433)),16);
when x"59a" => lut_sig <= to_unsigned(integer(my_cos(1434)),16);
when x"59b" => lut_sig <= to_unsigned(integer(my_cos(1435)),16);
when x"59c" => lut_sig <= to_unsigned(integer(my_cos(1436)),16);
when x"59d" => lut_sig <= to_unsigned(integer(my_cos(1437)),16);
when x"59e" => lut_sig <= to_unsigned(integer(my_cos(1438)),16);
when x"59f" => lut_sig <= to_unsigned(integer(my_cos(1439)),16);
when x"5a0" => lut_sig <= to_unsigned(integer(my_cos(1440)),16);
when x"5a1" => lut_sig <= to_unsigned(integer(my_cos(1441)),16);
when x"5a2" => lut_sig <= to_unsigned(integer(my_cos(1442)),16);
when x"5a3" => lut_sig <= to_unsigned(integer(my_cos(1443)),16);
when x"5a4" => lut_sig <= to_unsigned(integer(my_cos(1444)),16);
when x"5a5" => lut_sig <= to_unsigned(integer(my_cos(1445)),16);
when x"5a6" => lut_sig <= to_unsigned(integer(my_cos(1446)),16);
when x"5a7" => lut_sig <= to_unsigned(integer(my_cos(1447)),16);
when x"5a8" => lut_sig <= to_unsigned(integer(my_cos(1448)),16);
when x"5a9" => lut_sig <= to_unsigned(integer(my_cos(1449)),16);
when x"5aa" => lut_sig <= to_unsigned(integer(my_cos(1450)),16);
when x"5ab" => lut_sig <= to_unsigned(integer(my_cos(1451)),16);
when x"5ac" => lut_sig <= to_unsigned(integer(my_cos(1452)),16);
when x"5ad" => lut_sig <= to_unsigned(integer(my_cos(1453)),16);
when x"5ae" => lut_sig <= to_unsigned(integer(my_cos(1454)),16);
when x"5af" => lut_sig <= to_unsigned(integer(my_cos(1455)),16);
when x"5b0" => lut_sig <= to_unsigned(integer(my_cos(1456)),16);
when x"5b1" => lut_sig <= to_unsigned(integer(my_cos(1457)),16);
when x"5b2" => lut_sig <= to_unsigned(integer(my_cos(1458)),16);
when x"5b3" => lut_sig <= to_unsigned(integer(my_cos(1459)),16);
when x"5b4" => lut_sig <= to_unsigned(integer(my_cos(1460)),16);
when x"5b5" => lut_sig <= to_unsigned(integer(my_cos(1461)),16);
when x"5b6" => lut_sig <= to_unsigned(integer(my_cos(1462)),16);
when x"5b7" => lut_sig <= to_unsigned(integer(my_cos(1463)),16);
when x"5b8" => lut_sig <= to_unsigned(integer(my_cos(1464)),16);
when x"5b9" => lut_sig <= to_unsigned(integer(my_cos(1465)),16);
when x"5ba" => lut_sig <= to_unsigned(integer(my_cos(1466)),16);
when x"5bb" => lut_sig <= to_unsigned(integer(my_cos(1467)),16);
when x"5bc" => lut_sig <= to_unsigned(integer(my_cos(1468)),16);
when x"5bd" => lut_sig <= to_unsigned(integer(my_cos(1469)),16);
when x"5be" => lut_sig <= to_unsigned(integer(my_cos(1470)),16);
when x"5bf" => lut_sig <= to_unsigned(integer(my_cos(1471)),16);
when x"5c0" => lut_sig <= to_unsigned(integer(my_cos(1472)),16);
when x"5c1" => lut_sig <= to_unsigned(integer(my_cos(1473)),16);
when x"5c2" => lut_sig <= to_unsigned(integer(my_cos(1474)),16);
when x"5c3" => lut_sig <= to_unsigned(integer(my_cos(1475)),16);
when x"5c4" => lut_sig <= to_unsigned(integer(my_cos(1476)),16);
when x"5c5" => lut_sig <= to_unsigned(integer(my_cos(1477)),16);
when x"5c6" => lut_sig <= to_unsigned(integer(my_cos(1478)),16);
when x"5c7" => lut_sig <= to_unsigned(integer(my_cos(1479)),16);
when x"5c8" => lut_sig <= to_unsigned(integer(my_cos(1480)),16);
when x"5c9" => lut_sig <= to_unsigned(integer(my_cos(1481)),16);
when x"5ca" => lut_sig <= to_unsigned(integer(my_cos(1482)),16);
when x"5cb" => lut_sig <= to_unsigned(integer(my_cos(1483)),16);
when x"5cc" => lut_sig <= to_unsigned(integer(my_cos(1484)),16);
when x"5cd" => lut_sig <= to_unsigned(integer(my_cos(1485)),16);
when x"5ce" => lut_sig <= to_unsigned(integer(my_cos(1486)),16);
when x"5cf" => lut_sig <= to_unsigned(integer(my_cos(1487)),16);
when x"5d0" => lut_sig <= to_unsigned(integer(my_cos(1488)),16);
when x"5d1" => lut_sig <= to_unsigned(integer(my_cos(1489)),16);
when x"5d2" => lut_sig <= to_unsigned(integer(my_cos(1490)),16);
when x"5d3" => lut_sig <= to_unsigned(integer(my_cos(1491)),16);
when x"5d4" => lut_sig <= to_unsigned(integer(my_cos(1492)),16);
when x"5d5" => lut_sig <= to_unsigned(integer(my_cos(1493)),16);
when x"5d6" => lut_sig <= to_unsigned(integer(my_cos(1494)),16);
when x"5d7" => lut_sig <= to_unsigned(integer(my_cos(1495)),16);
when x"5d8" => lut_sig <= to_unsigned(integer(my_cos(1496)),16);
when x"5d9" => lut_sig <= to_unsigned(integer(my_cos(1497)),16);
when x"5da" => lut_sig <= to_unsigned(integer(my_cos(1498)),16);
when x"5db" => lut_sig <= to_unsigned(integer(my_cos(1499)),16);
when x"5dc" => lut_sig <= to_unsigned(integer(my_cos(1500)),16);
when x"5dd" => lut_sig <= to_unsigned(integer(my_cos(1501)),16);
when x"5de" => lut_sig <= to_unsigned(integer(my_cos(1502)),16);
when x"5df" => lut_sig <= to_unsigned(integer(my_cos(1503)),16);
when x"5e0" => lut_sig <= to_unsigned(integer(my_cos(1504)),16);
when x"5e1" => lut_sig <= to_unsigned(integer(my_cos(1505)),16);
when x"5e2" => lut_sig <= to_unsigned(integer(my_cos(1506)),16);
when x"5e3" => lut_sig <= to_unsigned(integer(my_cos(1507)),16);
when x"5e4" => lut_sig <= to_unsigned(integer(my_cos(1508)),16);
when x"5e5" => lut_sig <= to_unsigned(integer(my_cos(1509)),16);
when x"5e6" => lut_sig <= to_unsigned(integer(my_cos(1510)),16);
when x"5e7" => lut_sig <= to_unsigned(integer(my_cos(1511)),16);
when x"5e8" => lut_sig <= to_unsigned(integer(my_cos(1512)),16);
when x"5e9" => lut_sig <= to_unsigned(integer(my_cos(1513)),16);
when x"5ea" => lut_sig <= to_unsigned(integer(my_cos(1514)),16);
when x"5eb" => lut_sig <= to_unsigned(integer(my_cos(1515)),16);
when x"5ec" => lut_sig <= to_unsigned(integer(my_cos(1516)),16);
when x"5ed" => lut_sig <= to_unsigned(integer(my_cos(1517)),16);
when x"5ee" => lut_sig <= to_unsigned(integer(my_cos(1518)),16);
when x"5ef" => lut_sig <= to_unsigned(integer(my_cos(1519)),16);
when x"5f0" => lut_sig <= to_unsigned(integer(my_cos(1520)),16);
when x"5f1" => lut_sig <= to_unsigned(integer(my_cos(1521)),16);
when x"5f2" => lut_sig <= to_unsigned(integer(my_cos(1522)),16);
when x"5f3" => lut_sig <= to_unsigned(integer(my_cos(1523)),16);
when x"5f4" => lut_sig <= to_unsigned(integer(my_cos(1524)),16);
when x"5f5" => lut_sig <= to_unsigned(integer(my_cos(1525)),16);
when x"5f6" => lut_sig <= to_unsigned(integer(my_cos(1526)),16);
when x"5f7" => lut_sig <= to_unsigned(integer(my_cos(1527)),16);
when x"5f8" => lut_sig <= to_unsigned(integer(my_cos(1528)),16);
when x"5f9" => lut_sig <= to_unsigned(integer(my_cos(1529)),16);
when x"5fa" => lut_sig <= to_unsigned(integer(my_cos(1530)),16);
when x"5fb" => lut_sig <= to_unsigned(integer(my_cos(1531)),16);
when x"5fc" => lut_sig <= to_unsigned(integer(my_cos(1532)),16);
when x"5fd" => lut_sig <= to_unsigned(integer(my_cos(1533)),16);
when x"5fe" => lut_sig <= to_unsigned(integer(my_cos(1534)),16);
when x"5ff" => lut_sig <= to_unsigned(integer(my_cos(1535)),16);
when x"600" => lut_sig <= to_unsigned(integer(my_cos(1536)),16);
when x"601" => lut_sig <= to_unsigned(integer(my_cos(1537)),16);
when x"602" => lut_sig <= to_unsigned(integer(my_cos(1538)),16);
when x"603" => lut_sig <= to_unsigned(integer(my_cos(1539)),16);
when x"604" => lut_sig <= to_unsigned(integer(my_cos(1540)),16);
when x"605" => lut_sig <= to_unsigned(integer(my_cos(1541)),16);
when x"606" => lut_sig <= to_unsigned(integer(my_cos(1542)),16);
when x"607" => lut_sig <= to_unsigned(integer(my_cos(1543)),16);
when x"608" => lut_sig <= to_unsigned(integer(my_cos(1544)),16);
when x"609" => lut_sig <= to_unsigned(integer(my_cos(1545)),16);
when x"60a" => lut_sig <= to_unsigned(integer(my_cos(1546)),16);
when x"60b" => lut_sig <= to_unsigned(integer(my_cos(1547)),16);
when x"60c" => lut_sig <= to_unsigned(integer(my_cos(1548)),16);
when x"60d" => lut_sig <= to_unsigned(integer(my_cos(1549)),16);
when x"60e" => lut_sig <= to_unsigned(integer(my_cos(1550)),16);
when x"60f" => lut_sig <= to_unsigned(integer(my_cos(1551)),16);
when x"610" => lut_sig <= to_unsigned(integer(my_cos(1552)),16);
when x"611" => lut_sig <= to_unsigned(integer(my_cos(1553)),16);
when x"612" => lut_sig <= to_unsigned(integer(my_cos(1554)),16);
when x"613" => lut_sig <= to_unsigned(integer(my_cos(1555)),16);
when x"614" => lut_sig <= to_unsigned(integer(my_cos(1556)),16);
when x"615" => lut_sig <= to_unsigned(integer(my_cos(1557)),16);
when x"616" => lut_sig <= to_unsigned(integer(my_cos(1558)),16);
when x"617" => lut_sig <= to_unsigned(integer(my_cos(1559)),16);
when x"618" => lut_sig <= to_unsigned(integer(my_cos(1560)),16);
when x"619" => lut_sig <= to_unsigned(integer(my_cos(1561)),16);
when x"61a" => lut_sig <= to_unsigned(integer(my_cos(1562)),16);
when x"61b" => lut_sig <= to_unsigned(integer(my_cos(1563)),16);
when x"61c" => lut_sig <= to_unsigned(integer(my_cos(1564)),16);
when x"61d" => lut_sig <= to_unsigned(integer(my_cos(1565)),16);
when x"61e" => lut_sig <= to_unsigned(integer(my_cos(1566)),16);
when x"61f" => lut_sig <= to_unsigned(integer(my_cos(1567)),16);
when x"620" => lut_sig <= to_unsigned(integer(my_cos(1568)),16);
when x"621" => lut_sig <= to_unsigned(integer(my_cos(1569)),16);
when x"622" => lut_sig <= to_unsigned(integer(my_cos(1570)),16);
when x"623" => lut_sig <= to_unsigned(integer(my_cos(1571)),16);
when x"624" => lut_sig <= to_unsigned(integer(my_cos(1572)),16);
when x"625" => lut_sig <= to_unsigned(integer(my_cos(1573)),16);
when x"626" => lut_sig <= to_unsigned(integer(my_cos(1574)),16);
when x"627" => lut_sig <= to_unsigned(integer(my_cos(1575)),16);
when x"628" => lut_sig <= to_unsigned(integer(my_cos(1576)),16);
when x"629" => lut_sig <= to_unsigned(integer(my_cos(1577)),16);
when x"62a" => lut_sig <= to_unsigned(integer(my_cos(1578)),16);
when x"62b" => lut_sig <= to_unsigned(integer(my_cos(1579)),16);
when x"62c" => lut_sig <= to_unsigned(integer(my_cos(1580)),16);
when x"62d" => lut_sig <= to_unsigned(integer(my_cos(1581)),16);
when x"62e" => lut_sig <= to_unsigned(integer(my_cos(1582)),16);
when x"62f" => lut_sig <= to_unsigned(integer(my_cos(1583)),16);
when x"630" => lut_sig <= to_unsigned(integer(my_cos(1584)),16);
when x"631" => lut_sig <= to_unsigned(integer(my_cos(1585)),16);
when x"632" => lut_sig <= to_unsigned(integer(my_cos(1586)),16);
when x"633" => lut_sig <= to_unsigned(integer(my_cos(1587)),16);
when x"634" => lut_sig <= to_unsigned(integer(my_cos(1588)),16);
when x"635" => lut_sig <= to_unsigned(integer(my_cos(1589)),16);
when x"636" => lut_sig <= to_unsigned(integer(my_cos(1590)),16);
when x"637" => lut_sig <= to_unsigned(integer(my_cos(1591)),16);
when x"638" => lut_sig <= to_unsigned(integer(my_cos(1592)),16);
when x"639" => lut_sig <= to_unsigned(integer(my_cos(1593)),16);
when x"63a" => lut_sig <= to_unsigned(integer(my_cos(1594)),16);
when x"63b" => lut_sig <= to_unsigned(integer(my_cos(1595)),16);
when x"63c" => lut_sig <= to_unsigned(integer(my_cos(1596)),16);
when x"63d" => lut_sig <= to_unsigned(integer(my_cos(1597)),16);
when x"63e" => lut_sig <= to_unsigned(integer(my_cos(1598)),16);
when x"63f" => lut_sig <= to_unsigned(integer(my_cos(1599)),16);
when x"640" => lut_sig <= to_unsigned(integer(my_cos(1600)),16);
when x"641" => lut_sig <= to_unsigned(integer(my_cos(1601)),16);
when x"642" => lut_sig <= to_unsigned(integer(my_cos(1602)),16);
when x"643" => lut_sig <= to_unsigned(integer(my_cos(1603)),16);
when x"644" => lut_sig <= to_unsigned(integer(my_cos(1604)),16);
when x"645" => lut_sig <= to_unsigned(integer(my_cos(1605)),16);
when x"646" => lut_sig <= to_unsigned(integer(my_cos(1606)),16);
when x"647" => lut_sig <= to_unsigned(integer(my_cos(1607)),16);
when x"648" => lut_sig <= to_unsigned(integer(my_cos(1608)),16);
when x"649" => lut_sig <= to_unsigned(integer(my_cos(1609)),16);
when x"64a" => lut_sig <= to_unsigned(integer(my_cos(1610)),16);
when x"64b" => lut_sig <= to_unsigned(integer(my_cos(1611)),16);
when x"64c" => lut_sig <= to_unsigned(integer(my_cos(1612)),16);
when x"64d" => lut_sig <= to_unsigned(integer(my_cos(1613)),16);
when x"64e" => lut_sig <= to_unsigned(integer(my_cos(1614)),16);
when x"64f" => lut_sig <= to_unsigned(integer(my_cos(1615)),16);
when x"650" => lut_sig <= to_unsigned(integer(my_cos(1616)),16);
when x"651" => lut_sig <= to_unsigned(integer(my_cos(1617)),16);
when x"652" => lut_sig <= to_unsigned(integer(my_cos(1618)),16);
when x"653" => lut_sig <= to_unsigned(integer(my_cos(1619)),16);
when x"654" => lut_sig <= to_unsigned(integer(my_cos(1620)),16);
when x"655" => lut_sig <= to_unsigned(integer(my_cos(1621)),16);
when x"656" => lut_sig <= to_unsigned(integer(my_cos(1622)),16);
when x"657" => lut_sig <= to_unsigned(integer(my_cos(1623)),16);
when x"658" => lut_sig <= to_unsigned(integer(my_cos(1624)),16);
when x"659" => lut_sig <= to_unsigned(integer(my_cos(1625)),16);
when x"65a" => lut_sig <= to_unsigned(integer(my_cos(1626)),16);
when x"65b" => lut_sig <= to_unsigned(integer(my_cos(1627)),16);
when x"65c" => lut_sig <= to_unsigned(integer(my_cos(1628)),16);
when x"65d" => lut_sig <= to_unsigned(integer(my_cos(1629)),16);
when x"65e" => lut_sig <= to_unsigned(integer(my_cos(1630)),16);
when x"65f" => lut_sig <= to_unsigned(integer(my_cos(1631)),16);
when x"660" => lut_sig <= to_unsigned(integer(my_cos(1632)),16);
when x"661" => lut_sig <= to_unsigned(integer(my_cos(1633)),16);
when x"662" => lut_sig <= to_unsigned(integer(my_cos(1634)),16);
when x"663" => lut_sig <= to_unsigned(integer(my_cos(1635)),16);
when x"664" => lut_sig <= to_unsigned(integer(my_cos(1636)),16);
when x"665" => lut_sig <= to_unsigned(integer(my_cos(1637)),16);
when x"666" => lut_sig <= to_unsigned(integer(my_cos(1638)),16);
when x"667" => lut_sig <= to_unsigned(integer(my_cos(1639)),16);
when x"668" => lut_sig <= to_unsigned(integer(my_cos(1640)),16);
when x"669" => lut_sig <= to_unsigned(integer(my_cos(1641)),16);
when x"66a" => lut_sig <= to_unsigned(integer(my_cos(1642)),16);
when x"66b" => lut_sig <= to_unsigned(integer(my_cos(1643)),16);
when x"66c" => lut_sig <= to_unsigned(integer(my_cos(1644)),16);
when x"66d" => lut_sig <= to_unsigned(integer(my_cos(1645)),16);
when x"66e" => lut_sig <= to_unsigned(integer(my_cos(1646)),16);
when x"66f" => lut_sig <= to_unsigned(integer(my_cos(1647)),16);
when x"670" => lut_sig <= to_unsigned(integer(my_cos(1648)),16);
when x"671" => lut_sig <= to_unsigned(integer(my_cos(1649)),16);
when x"672" => lut_sig <= to_unsigned(integer(my_cos(1650)),16);
when x"673" => lut_sig <= to_unsigned(integer(my_cos(1651)),16);
when x"674" => lut_sig <= to_unsigned(integer(my_cos(1652)),16);
when x"675" => lut_sig <= to_unsigned(integer(my_cos(1653)),16);
when x"676" => lut_sig <= to_unsigned(integer(my_cos(1654)),16);
when x"677" => lut_sig <= to_unsigned(integer(my_cos(1655)),16);
when x"678" => lut_sig <= to_unsigned(integer(my_cos(1656)),16);
when x"679" => lut_sig <= to_unsigned(integer(my_cos(1657)),16);
when x"67a" => lut_sig <= to_unsigned(integer(my_cos(1658)),16);
when x"67b" => lut_sig <= to_unsigned(integer(my_cos(1659)),16);
when x"67c" => lut_sig <= to_unsigned(integer(my_cos(1660)),16);
when x"67d" => lut_sig <= to_unsigned(integer(my_cos(1661)),16);
when x"67e" => lut_sig <= to_unsigned(integer(my_cos(1662)),16);
when x"67f" => lut_sig <= to_unsigned(integer(my_cos(1663)),16);
when x"680" => lut_sig <= to_unsigned(integer(my_cos(1664)),16);
when x"681" => lut_sig <= to_unsigned(integer(my_cos(1665)),16);
when x"682" => lut_sig <= to_unsigned(integer(my_cos(1666)),16);
when x"683" => lut_sig <= to_unsigned(integer(my_cos(1667)),16);
when x"684" => lut_sig <= to_unsigned(integer(my_cos(1668)),16);
when x"685" => lut_sig <= to_unsigned(integer(my_cos(1669)),16);
when x"686" => lut_sig <= to_unsigned(integer(my_cos(1670)),16);
when x"687" => lut_sig <= to_unsigned(integer(my_cos(1671)),16);
when x"688" => lut_sig <= to_unsigned(integer(my_cos(1672)),16);
when x"689" => lut_sig <= to_unsigned(integer(my_cos(1673)),16);
when x"68a" => lut_sig <= to_unsigned(integer(my_cos(1674)),16);
when x"68b" => lut_sig <= to_unsigned(integer(my_cos(1675)),16);
when x"68c" => lut_sig <= to_unsigned(integer(my_cos(1676)),16);
when x"68d" => lut_sig <= to_unsigned(integer(my_cos(1677)),16);
when x"68e" => lut_sig <= to_unsigned(integer(my_cos(1678)),16);
when x"68f" => lut_sig <= to_unsigned(integer(my_cos(1679)),16);
when x"690" => lut_sig <= to_unsigned(integer(my_cos(1680)),16);
when x"691" => lut_sig <= to_unsigned(integer(my_cos(1681)),16);
when x"692" => lut_sig <= to_unsigned(integer(my_cos(1682)),16);
when x"693" => lut_sig <= to_unsigned(integer(my_cos(1683)),16);
when x"694" => lut_sig <= to_unsigned(integer(my_cos(1684)),16);
when x"695" => lut_sig <= to_unsigned(integer(my_cos(1685)),16);
when x"696" => lut_sig <= to_unsigned(integer(my_cos(1686)),16);
when x"697" => lut_sig <= to_unsigned(integer(my_cos(1687)),16);
when x"698" => lut_sig <= to_unsigned(integer(my_cos(1688)),16);
when x"699" => lut_sig <= to_unsigned(integer(my_cos(1689)),16);
when x"69a" => lut_sig <= to_unsigned(integer(my_cos(1690)),16);
when x"69b" => lut_sig <= to_unsigned(integer(my_cos(1691)),16);
when x"69c" => lut_sig <= to_unsigned(integer(my_cos(1692)),16);
when x"69d" => lut_sig <= to_unsigned(integer(my_cos(1693)),16);
when x"69e" => lut_sig <= to_unsigned(integer(my_cos(1694)),16);
when x"69f" => lut_sig <= to_unsigned(integer(my_cos(1695)),16);
when x"6a0" => lut_sig <= to_unsigned(integer(my_cos(1696)),16);
when x"6a1" => lut_sig <= to_unsigned(integer(my_cos(1697)),16);
when x"6a2" => lut_sig <= to_unsigned(integer(my_cos(1698)),16);
when x"6a3" => lut_sig <= to_unsigned(integer(my_cos(1699)),16);
when x"6a4" => lut_sig <= to_unsigned(integer(my_cos(1700)),16);
when x"6a5" => lut_sig <= to_unsigned(integer(my_cos(1701)),16);
when x"6a6" => lut_sig <= to_unsigned(integer(my_cos(1702)),16);
when x"6a7" => lut_sig <= to_unsigned(integer(my_cos(1703)),16);
when x"6a8" => lut_sig <= to_unsigned(integer(my_cos(1704)),16);
when x"6a9" => lut_sig <= to_unsigned(integer(my_cos(1705)),16);
when x"6aa" => lut_sig <= to_unsigned(integer(my_cos(1706)),16);
when x"6ab" => lut_sig <= to_unsigned(integer(my_cos(1707)),16);
when x"6ac" => lut_sig <= to_unsigned(integer(my_cos(1708)),16);
when x"6ad" => lut_sig <= to_unsigned(integer(my_cos(1709)),16);
when x"6ae" => lut_sig <= to_unsigned(integer(my_cos(1710)),16);
when x"6af" => lut_sig <= to_unsigned(integer(my_cos(1711)),16);
when x"6b0" => lut_sig <= to_unsigned(integer(my_cos(1712)),16);
when x"6b1" => lut_sig <= to_unsigned(integer(my_cos(1713)),16);
when x"6b2" => lut_sig <= to_unsigned(integer(my_cos(1714)),16);
when x"6b3" => lut_sig <= to_unsigned(integer(my_cos(1715)),16);
when x"6b4" => lut_sig <= to_unsigned(integer(my_cos(1716)),16);
when x"6b5" => lut_sig <= to_unsigned(integer(my_cos(1717)),16);
when x"6b6" => lut_sig <= to_unsigned(integer(my_cos(1718)),16);
when x"6b7" => lut_sig <= to_unsigned(integer(my_cos(1719)),16);
when x"6b8" => lut_sig <= to_unsigned(integer(my_cos(1720)),16);
when x"6b9" => lut_sig <= to_unsigned(integer(my_cos(1721)),16);
when x"6ba" => lut_sig <= to_unsigned(integer(my_cos(1722)),16);
when x"6bb" => lut_sig <= to_unsigned(integer(my_cos(1723)),16);
when x"6bc" => lut_sig <= to_unsigned(integer(my_cos(1724)),16);
when x"6bd" => lut_sig <= to_unsigned(integer(my_cos(1725)),16);
when x"6be" => lut_sig <= to_unsigned(integer(my_cos(1726)),16);
when x"6bf" => lut_sig <= to_unsigned(integer(my_cos(1727)),16);
when x"6c0" => lut_sig <= to_unsigned(integer(my_cos(1728)),16);
when x"6c1" => lut_sig <= to_unsigned(integer(my_cos(1729)),16);
when x"6c2" => lut_sig <= to_unsigned(integer(my_cos(1730)),16);
when x"6c3" => lut_sig <= to_unsigned(integer(my_cos(1731)),16);
when x"6c4" => lut_sig <= to_unsigned(integer(my_cos(1732)),16);
when x"6c5" => lut_sig <= to_unsigned(integer(my_cos(1733)),16);
when x"6c6" => lut_sig <= to_unsigned(integer(my_cos(1734)),16);
when x"6c7" => lut_sig <= to_unsigned(integer(my_cos(1735)),16);
when x"6c8" => lut_sig <= to_unsigned(integer(my_cos(1736)),16);
when x"6c9" => lut_sig <= to_unsigned(integer(my_cos(1737)),16);
when x"6ca" => lut_sig <= to_unsigned(integer(my_cos(1738)),16);
when x"6cb" => lut_sig <= to_unsigned(integer(my_cos(1739)),16);
when x"6cc" => lut_sig <= to_unsigned(integer(my_cos(1740)),16);
when x"6cd" => lut_sig <= to_unsigned(integer(my_cos(1741)),16);
when x"6ce" => lut_sig <= to_unsigned(integer(my_cos(1742)),16);
when x"6cf" => lut_sig <= to_unsigned(integer(my_cos(1743)),16);
when x"6d0" => lut_sig <= to_unsigned(integer(my_cos(1744)),16);
when x"6d1" => lut_sig <= to_unsigned(integer(my_cos(1745)),16);
when x"6d2" => lut_sig <= to_unsigned(integer(my_cos(1746)),16);
when x"6d3" => lut_sig <= to_unsigned(integer(my_cos(1747)),16);
when x"6d4" => lut_sig <= to_unsigned(integer(my_cos(1748)),16);
when x"6d5" => lut_sig <= to_unsigned(integer(my_cos(1749)),16);
when x"6d6" => lut_sig <= to_unsigned(integer(my_cos(1750)),16);
when x"6d7" => lut_sig <= to_unsigned(integer(my_cos(1751)),16);
when x"6d8" => lut_sig <= to_unsigned(integer(my_cos(1752)),16);
when x"6d9" => lut_sig <= to_unsigned(integer(my_cos(1753)),16);
when x"6da" => lut_sig <= to_unsigned(integer(my_cos(1754)),16);
when x"6db" => lut_sig <= to_unsigned(integer(my_cos(1755)),16);
when x"6dc" => lut_sig <= to_unsigned(integer(my_cos(1756)),16);
when x"6dd" => lut_sig <= to_unsigned(integer(my_cos(1757)),16);
when x"6de" => lut_sig <= to_unsigned(integer(my_cos(1758)),16);
when x"6df" => lut_sig <= to_unsigned(integer(my_cos(1759)),16);
when x"6e0" => lut_sig <= to_unsigned(integer(my_cos(1760)),16);
when x"6e1" => lut_sig <= to_unsigned(integer(my_cos(1761)),16);
when x"6e2" => lut_sig <= to_unsigned(integer(my_cos(1762)),16);
when x"6e3" => lut_sig <= to_unsigned(integer(my_cos(1763)),16);
when x"6e4" => lut_sig <= to_unsigned(integer(my_cos(1764)),16);
when x"6e5" => lut_sig <= to_unsigned(integer(my_cos(1765)),16);
when x"6e6" => lut_sig <= to_unsigned(integer(my_cos(1766)),16);
when x"6e7" => lut_sig <= to_unsigned(integer(my_cos(1767)),16);
when x"6e8" => lut_sig <= to_unsigned(integer(my_cos(1768)),16);
when x"6e9" => lut_sig <= to_unsigned(integer(my_cos(1769)),16);
when x"6ea" => lut_sig <= to_unsigned(integer(my_cos(1770)),16);
when x"6eb" => lut_sig <= to_unsigned(integer(my_cos(1771)),16);
when x"6ec" => lut_sig <= to_unsigned(integer(my_cos(1772)),16);
when x"6ed" => lut_sig <= to_unsigned(integer(my_cos(1773)),16);
when x"6ee" => lut_sig <= to_unsigned(integer(my_cos(1774)),16);
when x"6ef" => lut_sig <= to_unsigned(integer(my_cos(1775)),16);
when x"6f0" => lut_sig <= to_unsigned(integer(my_cos(1776)),16);
when x"6f1" => lut_sig <= to_unsigned(integer(my_cos(1777)),16);
when x"6f2" => lut_sig <= to_unsigned(integer(my_cos(1778)),16);
when x"6f3" => lut_sig <= to_unsigned(integer(my_cos(1779)),16);
when x"6f4" => lut_sig <= to_unsigned(integer(my_cos(1780)),16);
when x"6f5" => lut_sig <= to_unsigned(integer(my_cos(1781)),16);
when x"6f6" => lut_sig <= to_unsigned(integer(my_cos(1782)),16);
when x"6f7" => lut_sig <= to_unsigned(integer(my_cos(1783)),16);
when x"6f8" => lut_sig <= to_unsigned(integer(my_cos(1784)),16);
when x"6f9" => lut_sig <= to_unsigned(integer(my_cos(1785)),16);
when x"6fa" => lut_sig <= to_unsigned(integer(my_cos(1786)),16);
when x"6fb" => lut_sig <= to_unsigned(integer(my_cos(1787)),16);
when x"6fc" => lut_sig <= to_unsigned(integer(my_cos(1788)),16);
when x"6fd" => lut_sig <= to_unsigned(integer(my_cos(1789)),16);
when x"6fe" => lut_sig <= to_unsigned(integer(my_cos(1790)),16);
when x"6ff" => lut_sig <= to_unsigned(integer(my_cos(1791)),16);
when x"700" => lut_sig <= to_unsigned(integer(my_cos(1792)),16);
when x"701" => lut_sig <= to_unsigned(integer(my_cos(1793)),16);
when x"702" => lut_sig <= to_unsigned(integer(my_cos(1794)),16);
when x"703" => lut_sig <= to_unsigned(integer(my_cos(1795)),16);
when x"704" => lut_sig <= to_unsigned(integer(my_cos(1796)),16);
when x"705" => lut_sig <= to_unsigned(integer(my_cos(1797)),16);
when x"706" => lut_sig <= to_unsigned(integer(my_cos(1798)),16);
when x"707" => lut_sig <= to_unsigned(integer(my_cos(1799)),16);
when x"708" => lut_sig <= to_unsigned(integer(my_cos(1800)),16);
when x"709" => lut_sig <= to_unsigned(integer(my_cos(1801)),16);
when x"70a" => lut_sig <= to_unsigned(integer(my_cos(1802)),16);
when x"70b" => lut_sig <= to_unsigned(integer(my_cos(1803)),16);
when x"70c" => lut_sig <= to_unsigned(integer(my_cos(1804)),16);
when x"70d" => lut_sig <= to_unsigned(integer(my_cos(1805)),16);
when x"70e" => lut_sig <= to_unsigned(integer(my_cos(1806)),16);
when x"70f" => lut_sig <= to_unsigned(integer(my_cos(1807)),16);
when x"710" => lut_sig <= to_unsigned(integer(my_cos(1808)),16);
when x"711" => lut_sig <= to_unsigned(integer(my_cos(1809)),16);
when x"712" => lut_sig <= to_unsigned(integer(my_cos(1810)),16);
when x"713" => lut_sig <= to_unsigned(integer(my_cos(1811)),16);
when x"714" => lut_sig <= to_unsigned(integer(my_cos(1812)),16);
when x"715" => lut_sig <= to_unsigned(integer(my_cos(1813)),16);
when x"716" => lut_sig <= to_unsigned(integer(my_cos(1814)),16);
when x"717" => lut_sig <= to_unsigned(integer(my_cos(1815)),16);
when x"718" => lut_sig <= to_unsigned(integer(my_cos(1816)),16);
when x"719" => lut_sig <= to_unsigned(integer(my_cos(1817)),16);
when x"71a" => lut_sig <= to_unsigned(integer(my_cos(1818)),16);
when x"71b" => lut_sig <= to_unsigned(integer(my_cos(1819)),16);
when x"71c" => lut_sig <= to_unsigned(integer(my_cos(1820)),16);
when x"71d" => lut_sig <= to_unsigned(integer(my_cos(1821)),16);
when x"71e" => lut_sig <= to_unsigned(integer(my_cos(1822)),16);
when x"71f" => lut_sig <= to_unsigned(integer(my_cos(1823)),16);
when x"720" => lut_sig <= to_unsigned(integer(my_cos(1824)),16);
when x"721" => lut_sig <= to_unsigned(integer(my_cos(1825)),16);
when x"722" => lut_sig <= to_unsigned(integer(my_cos(1826)),16);
when x"723" => lut_sig <= to_unsigned(integer(my_cos(1827)),16);
when x"724" => lut_sig <= to_unsigned(integer(my_cos(1828)),16);
when x"725" => lut_sig <= to_unsigned(integer(my_cos(1829)),16);
when x"726" => lut_sig <= to_unsigned(integer(my_cos(1830)),16);
when x"727" => lut_sig <= to_unsigned(integer(my_cos(1831)),16);
when x"728" => lut_sig <= to_unsigned(integer(my_cos(1832)),16);
when x"729" => lut_sig <= to_unsigned(integer(my_cos(1833)),16);
when x"72a" => lut_sig <= to_unsigned(integer(my_cos(1834)),16);
when x"72b" => lut_sig <= to_unsigned(integer(my_cos(1835)),16);
when x"72c" => lut_sig <= to_unsigned(integer(my_cos(1836)),16);
when x"72d" => lut_sig <= to_unsigned(integer(my_cos(1837)),16);
when x"72e" => lut_sig <= to_unsigned(integer(my_cos(1838)),16);
when x"72f" => lut_sig <= to_unsigned(integer(my_cos(1839)),16);
when x"730" => lut_sig <= to_unsigned(integer(my_cos(1840)),16);
when x"731" => lut_sig <= to_unsigned(integer(my_cos(1841)),16);
when x"732" => lut_sig <= to_unsigned(integer(my_cos(1842)),16);
when x"733" => lut_sig <= to_unsigned(integer(my_cos(1843)),16);
when x"734" => lut_sig <= to_unsigned(integer(my_cos(1844)),16);
when x"735" => lut_sig <= to_unsigned(integer(my_cos(1845)),16);
when x"736" => lut_sig <= to_unsigned(integer(my_cos(1846)),16);
when x"737" => lut_sig <= to_unsigned(integer(my_cos(1847)),16);
when x"738" => lut_sig <= to_unsigned(integer(my_cos(1848)),16);
when x"739" => lut_sig <= to_unsigned(integer(my_cos(1849)),16);
when x"73a" => lut_sig <= to_unsigned(integer(my_cos(1850)),16);
when x"73b" => lut_sig <= to_unsigned(integer(my_cos(1851)),16);
when x"73c" => lut_sig <= to_unsigned(integer(my_cos(1852)),16);
when x"73d" => lut_sig <= to_unsigned(integer(my_cos(1853)),16);
when x"73e" => lut_sig <= to_unsigned(integer(my_cos(1854)),16);
when x"73f" => lut_sig <= to_unsigned(integer(my_cos(1855)),16);
when x"740" => lut_sig <= to_unsigned(integer(my_cos(1856)),16);
when x"741" => lut_sig <= to_unsigned(integer(my_cos(1857)),16);
when x"742" => lut_sig <= to_unsigned(integer(my_cos(1858)),16);
when x"743" => lut_sig <= to_unsigned(integer(my_cos(1859)),16);
when x"744" => lut_sig <= to_unsigned(integer(my_cos(1860)),16);
when x"745" => lut_sig <= to_unsigned(integer(my_cos(1861)),16);
when x"746" => lut_sig <= to_unsigned(integer(my_cos(1862)),16);
when x"747" => lut_sig <= to_unsigned(integer(my_cos(1863)),16);
when x"748" => lut_sig <= to_unsigned(integer(my_cos(1864)),16);
when x"749" => lut_sig <= to_unsigned(integer(my_cos(1865)),16);
when x"74a" => lut_sig <= to_unsigned(integer(my_cos(1866)),16);
when x"74b" => lut_sig <= to_unsigned(integer(my_cos(1867)),16);
when x"74c" => lut_sig <= to_unsigned(integer(my_cos(1868)),16);
when x"74d" => lut_sig <= to_unsigned(integer(my_cos(1869)),16);
when x"74e" => lut_sig <= to_unsigned(integer(my_cos(1870)),16);
when x"74f" => lut_sig <= to_unsigned(integer(my_cos(1871)),16);
when x"750" => lut_sig <= to_unsigned(integer(my_cos(1872)),16);
when x"751" => lut_sig <= to_unsigned(integer(my_cos(1873)),16);
when x"752" => lut_sig <= to_unsigned(integer(my_cos(1874)),16);
when x"753" => lut_sig <= to_unsigned(integer(my_cos(1875)),16);
when x"754" => lut_sig <= to_unsigned(integer(my_cos(1876)),16);
when x"755" => lut_sig <= to_unsigned(integer(my_cos(1877)),16);
when x"756" => lut_sig <= to_unsigned(integer(my_cos(1878)),16);
when x"757" => lut_sig <= to_unsigned(integer(my_cos(1879)),16);
when x"758" => lut_sig <= to_unsigned(integer(my_cos(1880)),16);
when x"759" => lut_sig <= to_unsigned(integer(my_cos(1881)),16);
when x"75a" => lut_sig <= to_unsigned(integer(my_cos(1882)),16);
when x"75b" => lut_sig <= to_unsigned(integer(my_cos(1883)),16);
when x"75c" => lut_sig <= to_unsigned(integer(my_cos(1884)),16);
when x"75d" => lut_sig <= to_unsigned(integer(my_cos(1885)),16);
when x"75e" => lut_sig <= to_unsigned(integer(my_cos(1886)),16);
when x"75f" => lut_sig <= to_unsigned(integer(my_cos(1887)),16);
when x"760" => lut_sig <= to_unsigned(integer(my_cos(1888)),16);
when x"761" => lut_sig <= to_unsigned(integer(my_cos(1889)),16);
when x"762" => lut_sig <= to_unsigned(integer(my_cos(1890)),16);
when x"763" => lut_sig <= to_unsigned(integer(my_cos(1891)),16);
when x"764" => lut_sig <= to_unsigned(integer(my_cos(1892)),16);
when x"765" => lut_sig <= to_unsigned(integer(my_cos(1893)),16);
when x"766" => lut_sig <= to_unsigned(integer(my_cos(1894)),16);
when x"767" => lut_sig <= to_unsigned(integer(my_cos(1895)),16);
when x"768" => lut_sig <= to_unsigned(integer(my_cos(1896)),16);
when x"769" => lut_sig <= to_unsigned(integer(my_cos(1897)),16);
when x"76a" => lut_sig <= to_unsigned(integer(my_cos(1898)),16);
when x"76b" => lut_sig <= to_unsigned(integer(my_cos(1899)),16);
when x"76c" => lut_sig <= to_unsigned(integer(my_cos(1900)),16);
when x"76d" => lut_sig <= to_unsigned(integer(my_cos(1901)),16);
when x"76e" => lut_sig <= to_unsigned(integer(my_cos(1902)),16);
when x"76f" => lut_sig <= to_unsigned(integer(my_cos(1903)),16);
when x"770" => lut_sig <= to_unsigned(integer(my_cos(1904)),16);
when x"771" => lut_sig <= to_unsigned(integer(my_cos(1905)),16);
when x"772" => lut_sig <= to_unsigned(integer(my_cos(1906)),16);
when x"773" => lut_sig <= to_unsigned(integer(my_cos(1907)),16);
when x"774" => lut_sig <= to_unsigned(integer(my_cos(1908)),16);
when x"775" => lut_sig <= to_unsigned(integer(my_cos(1909)),16);
when x"776" => lut_sig <= to_unsigned(integer(my_cos(1910)),16);
when x"777" => lut_sig <= to_unsigned(integer(my_cos(1911)),16);
when x"778" => lut_sig <= to_unsigned(integer(my_cos(1912)),16);
when x"779" => lut_sig <= to_unsigned(integer(my_cos(1913)),16);
when x"77a" => lut_sig <= to_unsigned(integer(my_cos(1914)),16);
when x"77b" => lut_sig <= to_unsigned(integer(my_cos(1915)),16);
when x"77c" => lut_sig <= to_unsigned(integer(my_cos(1916)),16);
when x"77d" => lut_sig <= to_unsigned(integer(my_cos(1917)),16);
when x"77e" => lut_sig <= to_unsigned(integer(my_cos(1918)),16);
when x"77f" => lut_sig <= to_unsigned(integer(my_cos(1919)),16);
when x"780" => lut_sig <= to_unsigned(integer(my_cos(1920)),16);
when x"781" => lut_sig <= to_unsigned(integer(my_cos(1921)),16);
when x"782" => lut_sig <= to_unsigned(integer(my_cos(1922)),16);
when x"783" => lut_sig <= to_unsigned(integer(my_cos(1923)),16);
when x"784" => lut_sig <= to_unsigned(integer(my_cos(1924)),16);
when x"785" => lut_sig <= to_unsigned(integer(my_cos(1925)),16);
when x"786" => lut_sig <= to_unsigned(integer(my_cos(1926)),16);
when x"787" => lut_sig <= to_unsigned(integer(my_cos(1927)),16);
when x"788" => lut_sig <= to_unsigned(integer(my_cos(1928)),16);
when x"789" => lut_sig <= to_unsigned(integer(my_cos(1929)),16);
when x"78a" => lut_sig <= to_unsigned(integer(my_cos(1930)),16);
when x"78b" => lut_sig <= to_unsigned(integer(my_cos(1931)),16);
when x"78c" => lut_sig <= to_unsigned(integer(my_cos(1932)),16);
when x"78d" => lut_sig <= to_unsigned(integer(my_cos(1933)),16);
when x"78e" => lut_sig <= to_unsigned(integer(my_cos(1934)),16);
when x"78f" => lut_sig <= to_unsigned(integer(my_cos(1935)),16);
when x"790" => lut_sig <= to_unsigned(integer(my_cos(1936)),16);
when x"791" => lut_sig <= to_unsigned(integer(my_cos(1937)),16);
when x"792" => lut_sig <= to_unsigned(integer(my_cos(1938)),16);
when x"793" => lut_sig <= to_unsigned(integer(my_cos(1939)),16);
when x"794" => lut_sig <= to_unsigned(integer(my_cos(1940)),16);
when x"795" => lut_sig <= to_unsigned(integer(my_cos(1941)),16);
when x"796" => lut_sig <= to_unsigned(integer(my_cos(1942)),16);
when x"797" => lut_sig <= to_unsigned(integer(my_cos(1943)),16);
when x"798" => lut_sig <= to_unsigned(integer(my_cos(1944)),16);
when x"799" => lut_sig <= to_unsigned(integer(my_cos(1945)),16);
when x"79a" => lut_sig <= to_unsigned(integer(my_cos(1946)),16);
when x"79b" => lut_sig <= to_unsigned(integer(my_cos(1947)),16);
when x"79c" => lut_sig <= to_unsigned(integer(my_cos(1948)),16);
when x"79d" => lut_sig <= to_unsigned(integer(my_cos(1949)),16);
when x"79e" => lut_sig <= to_unsigned(integer(my_cos(1950)),16);
when x"79f" => lut_sig <= to_unsigned(integer(my_cos(1951)),16);
when x"7a0" => lut_sig <= to_unsigned(integer(my_cos(1952)),16);
when x"7a1" => lut_sig <= to_unsigned(integer(my_cos(1953)),16);
when x"7a2" => lut_sig <= to_unsigned(integer(my_cos(1954)),16);
when x"7a3" => lut_sig <= to_unsigned(integer(my_cos(1955)),16);
when x"7a4" => lut_sig <= to_unsigned(integer(my_cos(1956)),16);
when x"7a5" => lut_sig <= to_unsigned(integer(my_cos(1957)),16);
when x"7a6" => lut_sig <= to_unsigned(integer(my_cos(1958)),16);
when x"7a7" => lut_sig <= to_unsigned(integer(my_cos(1959)),16);
when x"7a8" => lut_sig <= to_unsigned(integer(my_cos(1960)),16);
when x"7a9" => lut_sig <= to_unsigned(integer(my_cos(1961)),16);
when x"7aa" => lut_sig <= to_unsigned(integer(my_cos(1962)),16);
when x"7ab" => lut_sig <= to_unsigned(integer(my_cos(1963)),16);
when x"7ac" => lut_sig <= to_unsigned(integer(my_cos(1964)),16);
when x"7ad" => lut_sig <= to_unsigned(integer(my_cos(1965)),16);
when x"7ae" => lut_sig <= to_unsigned(integer(my_cos(1966)),16);
when x"7af" => lut_sig <= to_unsigned(integer(my_cos(1967)),16);
when x"7b0" => lut_sig <= to_unsigned(integer(my_cos(1968)),16);
when x"7b1" => lut_sig <= to_unsigned(integer(my_cos(1969)),16);
when x"7b2" => lut_sig <= to_unsigned(integer(my_cos(1970)),16);
when x"7b3" => lut_sig <= to_unsigned(integer(my_cos(1971)),16);
when x"7b4" => lut_sig <= to_unsigned(integer(my_cos(1972)),16);
when x"7b5" => lut_sig <= to_unsigned(integer(my_cos(1973)),16);
when x"7b6" => lut_sig <= to_unsigned(integer(my_cos(1974)),16);
when x"7b7" => lut_sig <= to_unsigned(integer(my_cos(1975)),16);
when x"7b8" => lut_sig <= to_unsigned(integer(my_cos(1976)),16);
when x"7b9" => lut_sig <= to_unsigned(integer(my_cos(1977)),16);
when x"7ba" => lut_sig <= to_unsigned(integer(my_cos(1978)),16);
when x"7bb" => lut_sig <= to_unsigned(integer(my_cos(1979)),16);
when x"7bc" => lut_sig <= to_unsigned(integer(my_cos(1980)),16);
when x"7bd" => lut_sig <= to_unsigned(integer(my_cos(1981)),16);
when x"7be" => lut_sig <= to_unsigned(integer(my_cos(1982)),16);
when x"7bf" => lut_sig <= to_unsigned(integer(my_cos(1983)),16);
when x"7c0" => lut_sig <= to_unsigned(integer(my_cos(1984)),16);
when x"7c1" => lut_sig <= to_unsigned(integer(my_cos(1985)),16);
when x"7c2" => lut_sig <= to_unsigned(integer(my_cos(1986)),16);
when x"7c3" => lut_sig <= to_unsigned(integer(my_cos(1987)),16);
when x"7c4" => lut_sig <= to_unsigned(integer(my_cos(1988)),16);
when x"7c5" => lut_sig <= to_unsigned(integer(my_cos(1989)),16);
when x"7c6" => lut_sig <= to_unsigned(integer(my_cos(1990)),16);
when x"7c7" => lut_sig <= to_unsigned(integer(my_cos(1991)),16);
when x"7c8" => lut_sig <= to_unsigned(integer(my_cos(1992)),16);
when x"7c9" => lut_sig <= to_unsigned(integer(my_cos(1993)),16);
when x"7ca" => lut_sig <= to_unsigned(integer(my_cos(1994)),16);
when x"7cb" => lut_sig <= to_unsigned(integer(my_cos(1995)),16);
when x"7cc" => lut_sig <= to_unsigned(integer(my_cos(1996)),16);
when x"7cd" => lut_sig <= to_unsigned(integer(my_cos(1997)),16);
when x"7ce" => lut_sig <= to_unsigned(integer(my_cos(1998)),16);
when x"7cf" => lut_sig <= to_unsigned(integer(my_cos(1999)),16);
when x"7d0" => lut_sig <= to_unsigned(integer(my_cos(2000)),16);
when x"7d1" => lut_sig <= to_unsigned(integer(my_cos(2001)),16);
when x"7d2" => lut_sig <= to_unsigned(integer(my_cos(2002)),16);
when x"7d3" => lut_sig <= to_unsigned(integer(my_cos(2003)),16);
when x"7d4" => lut_sig <= to_unsigned(integer(my_cos(2004)),16);
when x"7d5" => lut_sig <= to_unsigned(integer(my_cos(2005)),16);
when x"7d6" => lut_sig <= to_unsigned(integer(my_cos(2006)),16);
when x"7d7" => lut_sig <= to_unsigned(integer(my_cos(2007)),16);
when x"7d8" => lut_sig <= to_unsigned(integer(my_cos(2008)),16);
when x"7d9" => lut_sig <= to_unsigned(integer(my_cos(2009)),16);
when x"7da" => lut_sig <= to_unsigned(integer(my_cos(2010)),16);
when x"7db" => lut_sig <= to_unsigned(integer(my_cos(2011)),16);
when x"7dc" => lut_sig <= to_unsigned(integer(my_cos(2012)),16);
when x"7dd" => lut_sig <= to_unsigned(integer(my_cos(2013)),16);
when x"7de" => lut_sig <= to_unsigned(integer(my_cos(2014)),16);
when x"7df" => lut_sig <= to_unsigned(integer(my_cos(2015)),16);
when x"7e0" => lut_sig <= to_unsigned(integer(my_cos(2016)),16);
when x"7e1" => lut_sig <= to_unsigned(integer(my_cos(2017)),16);
when x"7e2" => lut_sig <= to_unsigned(integer(my_cos(2018)),16);
when x"7e3" => lut_sig <= to_unsigned(integer(my_cos(2019)),16);
when x"7e4" => lut_sig <= to_unsigned(integer(my_cos(2020)),16);
when x"7e5" => lut_sig <= to_unsigned(integer(my_cos(2021)),16);
when x"7e6" => lut_sig <= to_unsigned(integer(my_cos(2022)),16);
when x"7e7" => lut_sig <= to_unsigned(integer(my_cos(2023)),16);
when x"7e8" => lut_sig <= to_unsigned(integer(my_cos(2024)),16);
when x"7e9" => lut_sig <= to_unsigned(integer(my_cos(2025)),16);
when x"7ea" => lut_sig <= to_unsigned(integer(my_cos(2026)),16);
when x"7eb" => lut_sig <= to_unsigned(integer(my_cos(2027)),16);
when x"7ec" => lut_sig <= to_unsigned(integer(my_cos(2028)),16);
when x"7ed" => lut_sig <= to_unsigned(integer(my_cos(2029)),16);
when x"7ee" => lut_sig <= to_unsigned(integer(my_cos(2030)),16);
when x"7ef" => lut_sig <= to_unsigned(integer(my_cos(2031)),16);
when x"7f0" => lut_sig <= to_unsigned(integer(my_cos(2032)),16);
when x"7f1" => lut_sig <= to_unsigned(integer(my_cos(2033)),16);
when x"7f2" => lut_sig <= to_unsigned(integer(my_cos(2034)),16);
when x"7f3" => lut_sig <= to_unsigned(integer(my_cos(2035)),16);
when x"7f4" => lut_sig <= to_unsigned(integer(my_cos(2036)),16);
when x"7f5" => lut_sig <= to_unsigned(integer(my_cos(2037)),16);
when x"7f6" => lut_sig <= to_unsigned(integer(my_cos(2038)),16);
when x"7f7" => lut_sig <= to_unsigned(integer(my_cos(2039)),16);
when x"7f8" => lut_sig <= to_unsigned(integer(my_cos(2040)),16);
when x"7f9" => lut_sig <= to_unsigned(integer(my_cos(2041)),16);
when x"7fa" => lut_sig <= to_unsigned(integer(my_cos(2042)),16);
when x"7fb" => lut_sig <= to_unsigned(integer(my_cos(2043)),16);
when x"7fc" => lut_sig <= to_unsigned(integer(my_cos(2044)),16);
when x"7fd" => lut_sig <= to_unsigned(integer(my_cos(2045)),16);
when x"7fe" => lut_sig <= to_unsigned(integer(my_cos(2046)),16);
when x"7ff" => lut_sig <= to_unsigned(integer(my_cos(2047)),16);
when x"800" => lut_sig <= to_unsigned(integer(my_cos(2048)),16);
when x"801" => lut_sig <= to_unsigned(integer(my_cos(2049)),16);
when x"802" => lut_sig <= to_unsigned(integer(my_cos(2050)),16);
when x"803" => lut_sig <= to_unsigned(integer(my_cos(2051)),16);
when x"804" => lut_sig <= to_unsigned(integer(my_cos(2052)),16);
when x"805" => lut_sig <= to_unsigned(integer(my_cos(2053)),16);
when x"806" => lut_sig <= to_unsigned(integer(my_cos(2054)),16);
when x"807" => lut_sig <= to_unsigned(integer(my_cos(2055)),16);
when x"808" => lut_sig <= to_unsigned(integer(my_cos(2056)),16);
when x"809" => lut_sig <= to_unsigned(integer(my_cos(2057)),16);
when x"80a" => lut_sig <= to_unsigned(integer(my_cos(2058)),16);
when x"80b" => lut_sig <= to_unsigned(integer(my_cos(2059)),16);
when x"80c" => lut_sig <= to_unsigned(integer(my_cos(2060)),16);
when x"80d" => lut_sig <= to_unsigned(integer(my_cos(2061)),16);
when x"80e" => lut_sig <= to_unsigned(integer(my_cos(2062)),16);
when x"80f" => lut_sig <= to_unsigned(integer(my_cos(2063)),16);
when x"810" => lut_sig <= to_unsigned(integer(my_cos(2064)),16);
when x"811" => lut_sig <= to_unsigned(integer(my_cos(2065)),16);
when x"812" => lut_sig <= to_unsigned(integer(my_cos(2066)),16);
when x"813" => lut_sig <= to_unsigned(integer(my_cos(2067)),16);
when x"814" => lut_sig <= to_unsigned(integer(my_cos(2068)),16);
when x"815" => lut_sig <= to_unsigned(integer(my_cos(2069)),16);
when x"816" => lut_sig <= to_unsigned(integer(my_cos(2070)),16);
when x"817" => lut_sig <= to_unsigned(integer(my_cos(2071)),16);
when x"818" => lut_sig <= to_unsigned(integer(my_cos(2072)),16);
when x"819" => lut_sig <= to_unsigned(integer(my_cos(2073)),16);
when x"81a" => lut_sig <= to_unsigned(integer(my_cos(2074)),16);
when x"81b" => lut_sig <= to_unsigned(integer(my_cos(2075)),16);
when x"81c" => lut_sig <= to_unsigned(integer(my_cos(2076)),16);
when x"81d" => lut_sig <= to_unsigned(integer(my_cos(2077)),16);
when x"81e" => lut_sig <= to_unsigned(integer(my_cos(2078)),16);
when x"81f" => lut_sig <= to_unsigned(integer(my_cos(2079)),16);
when x"820" => lut_sig <= to_unsigned(integer(my_cos(2080)),16);
when x"821" => lut_sig <= to_unsigned(integer(my_cos(2081)),16);
when x"822" => lut_sig <= to_unsigned(integer(my_cos(2082)),16);
when x"823" => lut_sig <= to_unsigned(integer(my_cos(2083)),16);
when x"824" => lut_sig <= to_unsigned(integer(my_cos(2084)),16);
when x"825" => lut_sig <= to_unsigned(integer(my_cos(2085)),16);
when x"826" => lut_sig <= to_unsigned(integer(my_cos(2086)),16);
when x"827" => lut_sig <= to_unsigned(integer(my_cos(2087)),16);
when x"828" => lut_sig <= to_unsigned(integer(my_cos(2088)),16);
when x"829" => lut_sig <= to_unsigned(integer(my_cos(2089)),16);
when x"82a" => lut_sig <= to_unsigned(integer(my_cos(2090)),16);
when x"82b" => lut_sig <= to_unsigned(integer(my_cos(2091)),16);
when x"82c" => lut_sig <= to_unsigned(integer(my_cos(2092)),16);
when x"82d" => lut_sig <= to_unsigned(integer(my_cos(2093)),16);
when x"82e" => lut_sig <= to_unsigned(integer(my_cos(2094)),16);
when x"82f" => lut_sig <= to_unsigned(integer(my_cos(2095)),16);
when x"830" => lut_sig <= to_unsigned(integer(my_cos(2096)),16);
when x"831" => lut_sig <= to_unsigned(integer(my_cos(2097)),16);
when x"832" => lut_sig <= to_unsigned(integer(my_cos(2098)),16);
when x"833" => lut_sig <= to_unsigned(integer(my_cos(2099)),16);
when x"834" => lut_sig <= to_unsigned(integer(my_cos(2100)),16);
when x"835" => lut_sig <= to_unsigned(integer(my_cos(2101)),16);
when x"836" => lut_sig <= to_unsigned(integer(my_cos(2102)),16);
when x"837" => lut_sig <= to_unsigned(integer(my_cos(2103)),16);
when x"838" => lut_sig <= to_unsigned(integer(my_cos(2104)),16);
when x"839" => lut_sig <= to_unsigned(integer(my_cos(2105)),16);
when x"83a" => lut_sig <= to_unsigned(integer(my_cos(2106)),16);
when x"83b" => lut_sig <= to_unsigned(integer(my_cos(2107)),16);
when x"83c" => lut_sig <= to_unsigned(integer(my_cos(2108)),16);
when x"83d" => lut_sig <= to_unsigned(integer(my_cos(2109)),16);
when x"83e" => lut_sig <= to_unsigned(integer(my_cos(2110)),16);
when x"83f" => lut_sig <= to_unsigned(integer(my_cos(2111)),16);
when x"840" => lut_sig <= to_unsigned(integer(my_cos(2112)),16);
when x"841" => lut_sig <= to_unsigned(integer(my_cos(2113)),16);
when x"842" => lut_sig <= to_unsigned(integer(my_cos(2114)),16);
when x"843" => lut_sig <= to_unsigned(integer(my_cos(2115)),16);
when x"844" => lut_sig <= to_unsigned(integer(my_cos(2116)),16);
when x"845" => lut_sig <= to_unsigned(integer(my_cos(2117)),16);
when x"846" => lut_sig <= to_unsigned(integer(my_cos(2118)),16);
when x"847" => lut_sig <= to_unsigned(integer(my_cos(2119)),16);
when x"848" => lut_sig <= to_unsigned(integer(my_cos(2120)),16);
when x"849" => lut_sig <= to_unsigned(integer(my_cos(2121)),16);
when x"84a" => lut_sig <= to_unsigned(integer(my_cos(2122)),16);
when x"84b" => lut_sig <= to_unsigned(integer(my_cos(2123)),16);
when x"84c" => lut_sig <= to_unsigned(integer(my_cos(2124)),16);
when x"84d" => lut_sig <= to_unsigned(integer(my_cos(2125)),16);
when x"84e" => lut_sig <= to_unsigned(integer(my_cos(2126)),16);
when x"84f" => lut_sig <= to_unsigned(integer(my_cos(2127)),16);
when x"850" => lut_sig <= to_unsigned(integer(my_cos(2128)),16);
when x"851" => lut_sig <= to_unsigned(integer(my_cos(2129)),16);
when x"852" => lut_sig <= to_unsigned(integer(my_cos(2130)),16);
when x"853" => lut_sig <= to_unsigned(integer(my_cos(2131)),16);
when x"854" => lut_sig <= to_unsigned(integer(my_cos(2132)),16);
when x"855" => lut_sig <= to_unsigned(integer(my_cos(2133)),16);
when x"856" => lut_sig <= to_unsigned(integer(my_cos(2134)),16);
when x"857" => lut_sig <= to_unsigned(integer(my_cos(2135)),16);
when x"858" => lut_sig <= to_unsigned(integer(my_cos(2136)),16);
when x"859" => lut_sig <= to_unsigned(integer(my_cos(2137)),16);
when x"85a" => lut_sig <= to_unsigned(integer(my_cos(2138)),16);
when x"85b" => lut_sig <= to_unsigned(integer(my_cos(2139)),16);
when x"85c" => lut_sig <= to_unsigned(integer(my_cos(2140)),16);
when x"85d" => lut_sig <= to_unsigned(integer(my_cos(2141)),16);
when x"85e" => lut_sig <= to_unsigned(integer(my_cos(2142)),16);
when x"85f" => lut_sig <= to_unsigned(integer(my_cos(2143)),16);
when x"860" => lut_sig <= to_unsigned(integer(my_cos(2144)),16);
when x"861" => lut_sig <= to_unsigned(integer(my_cos(2145)),16);
when x"862" => lut_sig <= to_unsigned(integer(my_cos(2146)),16);
when x"863" => lut_sig <= to_unsigned(integer(my_cos(2147)),16);
when x"864" => lut_sig <= to_unsigned(integer(my_cos(2148)),16);
when x"865" => lut_sig <= to_unsigned(integer(my_cos(2149)),16);
when x"866" => lut_sig <= to_unsigned(integer(my_cos(2150)),16);
when x"867" => lut_sig <= to_unsigned(integer(my_cos(2151)),16);
when x"868" => lut_sig <= to_unsigned(integer(my_cos(2152)),16);
when x"869" => lut_sig <= to_unsigned(integer(my_cos(2153)),16);
when x"86a" => lut_sig <= to_unsigned(integer(my_cos(2154)),16);
when x"86b" => lut_sig <= to_unsigned(integer(my_cos(2155)),16);
when x"86c" => lut_sig <= to_unsigned(integer(my_cos(2156)),16);
when x"86d" => lut_sig <= to_unsigned(integer(my_cos(2157)),16);
when x"86e" => lut_sig <= to_unsigned(integer(my_cos(2158)),16);
when x"86f" => lut_sig <= to_unsigned(integer(my_cos(2159)),16);
when x"870" => lut_sig <= to_unsigned(integer(my_cos(2160)),16);
when x"871" => lut_sig <= to_unsigned(integer(my_cos(2161)),16);
when x"872" => lut_sig <= to_unsigned(integer(my_cos(2162)),16);
when x"873" => lut_sig <= to_unsigned(integer(my_cos(2163)),16);
when x"874" => lut_sig <= to_unsigned(integer(my_cos(2164)),16);
when x"875" => lut_sig <= to_unsigned(integer(my_cos(2165)),16);
when x"876" => lut_sig <= to_unsigned(integer(my_cos(2166)),16);
when x"877" => lut_sig <= to_unsigned(integer(my_cos(2167)),16);
when x"878" => lut_sig <= to_unsigned(integer(my_cos(2168)),16);
when x"879" => lut_sig <= to_unsigned(integer(my_cos(2169)),16);
when x"87a" => lut_sig <= to_unsigned(integer(my_cos(2170)),16);
when x"87b" => lut_sig <= to_unsigned(integer(my_cos(2171)),16);
when x"87c" => lut_sig <= to_unsigned(integer(my_cos(2172)),16);
when x"87d" => lut_sig <= to_unsigned(integer(my_cos(2173)),16);
when x"87e" => lut_sig <= to_unsigned(integer(my_cos(2174)),16);
when x"87f" => lut_sig <= to_unsigned(integer(my_cos(2175)),16);
when x"880" => lut_sig <= to_unsigned(integer(my_cos(2176)),16);
when x"881" => lut_sig <= to_unsigned(integer(my_cos(2177)),16);
when x"882" => lut_sig <= to_unsigned(integer(my_cos(2178)),16);
when x"883" => lut_sig <= to_unsigned(integer(my_cos(2179)),16);
when x"884" => lut_sig <= to_unsigned(integer(my_cos(2180)),16);
when x"885" => lut_sig <= to_unsigned(integer(my_cos(2181)),16);
when x"886" => lut_sig <= to_unsigned(integer(my_cos(2182)),16);
when x"887" => lut_sig <= to_unsigned(integer(my_cos(2183)),16);
when x"888" => lut_sig <= to_unsigned(integer(my_cos(2184)),16);
when x"889" => lut_sig <= to_unsigned(integer(my_cos(2185)),16);
when x"88a" => lut_sig <= to_unsigned(integer(my_cos(2186)),16);
when x"88b" => lut_sig <= to_unsigned(integer(my_cos(2187)),16);
when x"88c" => lut_sig <= to_unsigned(integer(my_cos(2188)),16);
when x"88d" => lut_sig <= to_unsigned(integer(my_cos(2189)),16);
when x"88e" => lut_sig <= to_unsigned(integer(my_cos(2190)),16);
when x"88f" => lut_sig <= to_unsigned(integer(my_cos(2191)),16);
when x"890" => lut_sig <= to_unsigned(integer(my_cos(2192)),16);
when x"891" => lut_sig <= to_unsigned(integer(my_cos(2193)),16);
when x"892" => lut_sig <= to_unsigned(integer(my_cos(2194)),16);
when x"893" => lut_sig <= to_unsigned(integer(my_cos(2195)),16);
when x"894" => lut_sig <= to_unsigned(integer(my_cos(2196)),16);
when x"895" => lut_sig <= to_unsigned(integer(my_cos(2197)),16);
when x"896" => lut_sig <= to_unsigned(integer(my_cos(2198)),16);
when x"897" => lut_sig <= to_unsigned(integer(my_cos(2199)),16);
when x"898" => lut_sig <= to_unsigned(integer(my_cos(2200)),16);
when x"899" => lut_sig <= to_unsigned(integer(my_cos(2201)),16);
when x"89a" => lut_sig <= to_unsigned(integer(my_cos(2202)),16);
when x"89b" => lut_sig <= to_unsigned(integer(my_cos(2203)),16);
when x"89c" => lut_sig <= to_unsigned(integer(my_cos(2204)),16);
when x"89d" => lut_sig <= to_unsigned(integer(my_cos(2205)),16);
when x"89e" => lut_sig <= to_unsigned(integer(my_cos(2206)),16);
when x"89f" => lut_sig <= to_unsigned(integer(my_cos(2207)),16);
when x"8a0" => lut_sig <= to_unsigned(integer(my_cos(2208)),16);
when x"8a1" => lut_sig <= to_unsigned(integer(my_cos(2209)),16);
when x"8a2" => lut_sig <= to_unsigned(integer(my_cos(2210)),16);
when x"8a3" => lut_sig <= to_unsigned(integer(my_cos(2211)),16);
when x"8a4" => lut_sig <= to_unsigned(integer(my_cos(2212)),16);
when x"8a5" => lut_sig <= to_unsigned(integer(my_cos(2213)),16);
when x"8a6" => lut_sig <= to_unsigned(integer(my_cos(2214)),16);
when x"8a7" => lut_sig <= to_unsigned(integer(my_cos(2215)),16);
when x"8a8" => lut_sig <= to_unsigned(integer(my_cos(2216)),16);
when x"8a9" => lut_sig <= to_unsigned(integer(my_cos(2217)),16);
when x"8aa" => lut_sig <= to_unsigned(integer(my_cos(2218)),16);
when x"8ab" => lut_sig <= to_unsigned(integer(my_cos(2219)),16);
when x"8ac" => lut_sig <= to_unsigned(integer(my_cos(2220)),16);
when x"8ad" => lut_sig <= to_unsigned(integer(my_cos(2221)),16);
when x"8ae" => lut_sig <= to_unsigned(integer(my_cos(2222)),16);
when x"8af" => lut_sig <= to_unsigned(integer(my_cos(2223)),16);
when x"8b0" => lut_sig <= to_unsigned(integer(my_cos(2224)),16);
when x"8b1" => lut_sig <= to_unsigned(integer(my_cos(2225)),16);
when x"8b2" => lut_sig <= to_unsigned(integer(my_cos(2226)),16);
when x"8b3" => lut_sig <= to_unsigned(integer(my_cos(2227)),16);
when x"8b4" => lut_sig <= to_unsigned(integer(my_cos(2228)),16);
when x"8b5" => lut_sig <= to_unsigned(integer(my_cos(2229)),16);
when x"8b6" => lut_sig <= to_unsigned(integer(my_cos(2230)),16);
when x"8b7" => lut_sig <= to_unsigned(integer(my_cos(2231)),16);
when x"8b8" => lut_sig <= to_unsigned(integer(my_cos(2232)),16);
when x"8b9" => lut_sig <= to_unsigned(integer(my_cos(2233)),16);
when x"8ba" => lut_sig <= to_unsigned(integer(my_cos(2234)),16);
when x"8bb" => lut_sig <= to_unsigned(integer(my_cos(2235)),16);
when x"8bc" => lut_sig <= to_unsigned(integer(my_cos(2236)),16);
when x"8bd" => lut_sig <= to_unsigned(integer(my_cos(2237)),16);
when x"8be" => lut_sig <= to_unsigned(integer(my_cos(2238)),16);
when x"8bf" => lut_sig <= to_unsigned(integer(my_cos(2239)),16);
when x"8c0" => lut_sig <= to_unsigned(integer(my_cos(2240)),16);
when x"8c1" => lut_sig <= to_unsigned(integer(my_cos(2241)),16);
when x"8c2" => lut_sig <= to_unsigned(integer(my_cos(2242)),16);
when x"8c3" => lut_sig <= to_unsigned(integer(my_cos(2243)),16);
when x"8c4" => lut_sig <= to_unsigned(integer(my_cos(2244)),16);
when x"8c5" => lut_sig <= to_unsigned(integer(my_cos(2245)),16);
when x"8c6" => lut_sig <= to_unsigned(integer(my_cos(2246)),16);
when x"8c7" => lut_sig <= to_unsigned(integer(my_cos(2247)),16);
when x"8c8" => lut_sig <= to_unsigned(integer(my_cos(2248)),16);
when x"8c9" => lut_sig <= to_unsigned(integer(my_cos(2249)),16);
when x"8ca" => lut_sig <= to_unsigned(integer(my_cos(2250)),16);
when x"8cb" => lut_sig <= to_unsigned(integer(my_cos(2251)),16);
when x"8cc" => lut_sig <= to_unsigned(integer(my_cos(2252)),16);
when x"8cd" => lut_sig <= to_unsigned(integer(my_cos(2253)),16);
when x"8ce" => lut_sig <= to_unsigned(integer(my_cos(2254)),16);
when x"8cf" => lut_sig <= to_unsigned(integer(my_cos(2255)),16);
when x"8d0" => lut_sig <= to_unsigned(integer(my_cos(2256)),16);
when x"8d1" => lut_sig <= to_unsigned(integer(my_cos(2257)),16);
when x"8d2" => lut_sig <= to_unsigned(integer(my_cos(2258)),16);
when x"8d3" => lut_sig <= to_unsigned(integer(my_cos(2259)),16);
when x"8d4" => lut_sig <= to_unsigned(integer(my_cos(2260)),16);
when x"8d5" => lut_sig <= to_unsigned(integer(my_cos(2261)),16);
when x"8d6" => lut_sig <= to_unsigned(integer(my_cos(2262)),16);
when x"8d7" => lut_sig <= to_unsigned(integer(my_cos(2263)),16);
when x"8d8" => lut_sig <= to_unsigned(integer(my_cos(2264)),16);
when x"8d9" => lut_sig <= to_unsigned(integer(my_cos(2265)),16);
when x"8da" => lut_sig <= to_unsigned(integer(my_cos(2266)),16);
when x"8db" => lut_sig <= to_unsigned(integer(my_cos(2267)),16);
when x"8dc" => lut_sig <= to_unsigned(integer(my_cos(2268)),16);
when x"8dd" => lut_sig <= to_unsigned(integer(my_cos(2269)),16);
when x"8de" => lut_sig <= to_unsigned(integer(my_cos(2270)),16);
when x"8df" => lut_sig <= to_unsigned(integer(my_cos(2271)),16);
when x"8e0" => lut_sig <= to_unsigned(integer(my_cos(2272)),16);
when x"8e1" => lut_sig <= to_unsigned(integer(my_cos(2273)),16);
when x"8e2" => lut_sig <= to_unsigned(integer(my_cos(2274)),16);
when x"8e3" => lut_sig <= to_unsigned(integer(my_cos(2275)),16);
when x"8e4" => lut_sig <= to_unsigned(integer(my_cos(2276)),16);
when x"8e5" => lut_sig <= to_unsigned(integer(my_cos(2277)),16);
when x"8e6" => lut_sig <= to_unsigned(integer(my_cos(2278)),16);
when x"8e7" => lut_sig <= to_unsigned(integer(my_cos(2279)),16);
when x"8e8" => lut_sig <= to_unsigned(integer(my_cos(2280)),16);
when x"8e9" => lut_sig <= to_unsigned(integer(my_cos(2281)),16);
when x"8ea" => lut_sig <= to_unsigned(integer(my_cos(2282)),16);
when x"8eb" => lut_sig <= to_unsigned(integer(my_cos(2283)),16);
when x"8ec" => lut_sig <= to_unsigned(integer(my_cos(2284)),16);
when x"8ed" => lut_sig <= to_unsigned(integer(my_cos(2285)),16);
when x"8ee" => lut_sig <= to_unsigned(integer(my_cos(2286)),16);
when x"8ef" => lut_sig <= to_unsigned(integer(my_cos(2287)),16);
when x"8f0" => lut_sig <= to_unsigned(integer(my_cos(2288)),16);
when x"8f1" => lut_sig <= to_unsigned(integer(my_cos(2289)),16);
when x"8f2" => lut_sig <= to_unsigned(integer(my_cos(2290)),16);
when x"8f3" => lut_sig <= to_unsigned(integer(my_cos(2291)),16);
when x"8f4" => lut_sig <= to_unsigned(integer(my_cos(2292)),16);
when x"8f5" => lut_sig <= to_unsigned(integer(my_cos(2293)),16);
when x"8f6" => lut_sig <= to_unsigned(integer(my_cos(2294)),16);
when x"8f7" => lut_sig <= to_unsigned(integer(my_cos(2295)),16);
when x"8f8" => lut_sig <= to_unsigned(integer(my_cos(2296)),16);
when x"8f9" => lut_sig <= to_unsigned(integer(my_cos(2297)),16);
when x"8fa" => lut_sig <= to_unsigned(integer(my_cos(2298)),16);
when x"8fb" => lut_sig <= to_unsigned(integer(my_cos(2299)),16);
when x"8fc" => lut_sig <= to_unsigned(integer(my_cos(2300)),16);
when x"8fd" => lut_sig <= to_unsigned(integer(my_cos(2301)),16);
when x"8fe" => lut_sig <= to_unsigned(integer(my_cos(2302)),16);
when x"8ff" => lut_sig <= to_unsigned(integer(my_cos(2303)),16);
when x"900" => lut_sig <= to_unsigned(integer(my_cos(2304)),16);
when x"901" => lut_sig <= to_unsigned(integer(my_cos(2305)),16);
when x"902" => lut_sig <= to_unsigned(integer(my_cos(2306)),16);
when x"903" => lut_sig <= to_unsigned(integer(my_cos(2307)),16);
when x"904" => lut_sig <= to_unsigned(integer(my_cos(2308)),16);
when x"905" => lut_sig <= to_unsigned(integer(my_cos(2309)),16);
when x"906" => lut_sig <= to_unsigned(integer(my_cos(2310)),16);
when x"907" => lut_sig <= to_unsigned(integer(my_cos(2311)),16);
when x"908" => lut_sig <= to_unsigned(integer(my_cos(2312)),16);
when x"909" => lut_sig <= to_unsigned(integer(my_cos(2313)),16);
when x"90a" => lut_sig <= to_unsigned(integer(my_cos(2314)),16);
when x"90b" => lut_sig <= to_unsigned(integer(my_cos(2315)),16);
when x"90c" => lut_sig <= to_unsigned(integer(my_cos(2316)),16);
when x"90d" => lut_sig <= to_unsigned(integer(my_cos(2317)),16);
when x"90e" => lut_sig <= to_unsigned(integer(my_cos(2318)),16);
when x"90f" => lut_sig <= to_unsigned(integer(my_cos(2319)),16);
when x"910" => lut_sig <= to_unsigned(integer(my_cos(2320)),16);
when x"911" => lut_sig <= to_unsigned(integer(my_cos(2321)),16);
when x"912" => lut_sig <= to_unsigned(integer(my_cos(2322)),16);
when x"913" => lut_sig <= to_unsigned(integer(my_cos(2323)),16);
when x"914" => lut_sig <= to_unsigned(integer(my_cos(2324)),16);
when x"915" => lut_sig <= to_unsigned(integer(my_cos(2325)),16);
when x"916" => lut_sig <= to_unsigned(integer(my_cos(2326)),16);
when x"917" => lut_sig <= to_unsigned(integer(my_cos(2327)),16);
when x"918" => lut_sig <= to_unsigned(integer(my_cos(2328)),16);
when x"919" => lut_sig <= to_unsigned(integer(my_cos(2329)),16);
when x"91a" => lut_sig <= to_unsigned(integer(my_cos(2330)),16);
when x"91b" => lut_sig <= to_unsigned(integer(my_cos(2331)),16);
when x"91c" => lut_sig <= to_unsigned(integer(my_cos(2332)),16);
when x"91d" => lut_sig <= to_unsigned(integer(my_cos(2333)),16);
when x"91e" => lut_sig <= to_unsigned(integer(my_cos(2334)),16);
when x"91f" => lut_sig <= to_unsigned(integer(my_cos(2335)),16);
when x"920" => lut_sig <= to_unsigned(integer(my_cos(2336)),16);
when x"921" => lut_sig <= to_unsigned(integer(my_cos(2337)),16);
when x"922" => lut_sig <= to_unsigned(integer(my_cos(2338)),16);
when x"923" => lut_sig <= to_unsigned(integer(my_cos(2339)),16);
when x"924" => lut_sig <= to_unsigned(integer(my_cos(2340)),16);
when x"925" => lut_sig <= to_unsigned(integer(my_cos(2341)),16);
when x"926" => lut_sig <= to_unsigned(integer(my_cos(2342)),16);
when x"927" => lut_sig <= to_unsigned(integer(my_cos(2343)),16);
when x"928" => lut_sig <= to_unsigned(integer(my_cos(2344)),16);
when x"929" => lut_sig <= to_unsigned(integer(my_cos(2345)),16);
when x"92a" => lut_sig <= to_unsigned(integer(my_cos(2346)),16);
when x"92b" => lut_sig <= to_unsigned(integer(my_cos(2347)),16);
when x"92c" => lut_sig <= to_unsigned(integer(my_cos(2348)),16);
when x"92d" => lut_sig <= to_unsigned(integer(my_cos(2349)),16);
when x"92e" => lut_sig <= to_unsigned(integer(my_cos(2350)),16);
when x"92f" => lut_sig <= to_unsigned(integer(my_cos(2351)),16);
when x"930" => lut_sig <= to_unsigned(integer(my_cos(2352)),16);
when x"931" => lut_sig <= to_unsigned(integer(my_cos(2353)),16);
when x"932" => lut_sig <= to_unsigned(integer(my_cos(2354)),16);
when x"933" => lut_sig <= to_unsigned(integer(my_cos(2355)),16);
when x"934" => lut_sig <= to_unsigned(integer(my_cos(2356)),16);
when x"935" => lut_sig <= to_unsigned(integer(my_cos(2357)),16);
when x"936" => lut_sig <= to_unsigned(integer(my_cos(2358)),16);
when x"937" => lut_sig <= to_unsigned(integer(my_cos(2359)),16);
when x"938" => lut_sig <= to_unsigned(integer(my_cos(2360)),16);
when x"939" => lut_sig <= to_unsigned(integer(my_cos(2361)),16);
when x"93a" => lut_sig <= to_unsigned(integer(my_cos(2362)),16);
when x"93b" => lut_sig <= to_unsigned(integer(my_cos(2363)),16);
when x"93c" => lut_sig <= to_unsigned(integer(my_cos(2364)),16);
when x"93d" => lut_sig <= to_unsigned(integer(my_cos(2365)),16);
when x"93e" => lut_sig <= to_unsigned(integer(my_cos(2366)),16);
when x"93f" => lut_sig <= to_unsigned(integer(my_cos(2367)),16);
when x"940" => lut_sig <= to_unsigned(integer(my_cos(2368)),16);
when x"941" => lut_sig <= to_unsigned(integer(my_cos(2369)),16);
when x"942" => lut_sig <= to_unsigned(integer(my_cos(2370)),16);
when x"943" => lut_sig <= to_unsigned(integer(my_cos(2371)),16);
when x"944" => lut_sig <= to_unsigned(integer(my_cos(2372)),16);
when x"945" => lut_sig <= to_unsigned(integer(my_cos(2373)),16);
when x"946" => lut_sig <= to_unsigned(integer(my_cos(2374)),16);
when x"947" => lut_sig <= to_unsigned(integer(my_cos(2375)),16);
when x"948" => lut_sig <= to_unsigned(integer(my_cos(2376)),16);
when x"949" => lut_sig <= to_unsigned(integer(my_cos(2377)),16);
when x"94a" => lut_sig <= to_unsigned(integer(my_cos(2378)),16);
when x"94b" => lut_sig <= to_unsigned(integer(my_cos(2379)),16);
when x"94c" => lut_sig <= to_unsigned(integer(my_cos(2380)),16);
when x"94d" => lut_sig <= to_unsigned(integer(my_cos(2381)),16);
when x"94e" => lut_sig <= to_unsigned(integer(my_cos(2382)),16);
when x"94f" => lut_sig <= to_unsigned(integer(my_cos(2383)),16);
when x"950" => lut_sig <= to_unsigned(integer(my_cos(2384)),16);
when x"951" => lut_sig <= to_unsigned(integer(my_cos(2385)),16);
when x"952" => lut_sig <= to_unsigned(integer(my_cos(2386)),16);
when x"953" => lut_sig <= to_unsigned(integer(my_cos(2387)),16);
when x"954" => lut_sig <= to_unsigned(integer(my_cos(2388)),16);
when x"955" => lut_sig <= to_unsigned(integer(my_cos(2389)),16);
when x"956" => lut_sig <= to_unsigned(integer(my_cos(2390)),16);
when x"957" => lut_sig <= to_unsigned(integer(my_cos(2391)),16);
when x"958" => lut_sig <= to_unsigned(integer(my_cos(2392)),16);
when x"959" => lut_sig <= to_unsigned(integer(my_cos(2393)),16);
when x"95a" => lut_sig <= to_unsigned(integer(my_cos(2394)),16);
when x"95b" => lut_sig <= to_unsigned(integer(my_cos(2395)),16);
when x"95c" => lut_sig <= to_unsigned(integer(my_cos(2396)),16);
when x"95d" => lut_sig <= to_unsigned(integer(my_cos(2397)),16);
when x"95e" => lut_sig <= to_unsigned(integer(my_cos(2398)),16);
when x"95f" => lut_sig <= to_unsigned(integer(my_cos(2399)),16);
when x"960" => lut_sig <= to_unsigned(integer(my_cos(2400)),16);
when x"961" => lut_sig <= to_unsigned(integer(my_cos(2401)),16);
when x"962" => lut_sig <= to_unsigned(integer(my_cos(2402)),16);
when x"963" => lut_sig <= to_unsigned(integer(my_cos(2403)),16);
when x"964" => lut_sig <= to_unsigned(integer(my_cos(2404)),16);
when x"965" => lut_sig <= to_unsigned(integer(my_cos(2405)),16);
when x"966" => lut_sig <= to_unsigned(integer(my_cos(2406)),16);
when x"967" => lut_sig <= to_unsigned(integer(my_cos(2407)),16);
when x"968" => lut_sig <= to_unsigned(integer(my_cos(2408)),16);
when x"969" => lut_sig <= to_unsigned(integer(my_cos(2409)),16);
when x"96a" => lut_sig <= to_unsigned(integer(my_cos(2410)),16);
when x"96b" => lut_sig <= to_unsigned(integer(my_cos(2411)),16);
when x"96c" => lut_sig <= to_unsigned(integer(my_cos(2412)),16);
when x"96d" => lut_sig <= to_unsigned(integer(my_cos(2413)),16);
when x"96e" => lut_sig <= to_unsigned(integer(my_cos(2414)),16);
when x"96f" => lut_sig <= to_unsigned(integer(my_cos(2415)),16);
when x"970" => lut_sig <= to_unsigned(integer(my_cos(2416)),16);
when x"971" => lut_sig <= to_unsigned(integer(my_cos(2417)),16);
when x"972" => lut_sig <= to_unsigned(integer(my_cos(2418)),16);
when x"973" => lut_sig <= to_unsigned(integer(my_cos(2419)),16);
when x"974" => lut_sig <= to_unsigned(integer(my_cos(2420)),16);
when x"975" => lut_sig <= to_unsigned(integer(my_cos(2421)),16);
when x"976" => lut_sig <= to_unsigned(integer(my_cos(2422)),16);
when x"977" => lut_sig <= to_unsigned(integer(my_cos(2423)),16);
when x"978" => lut_sig <= to_unsigned(integer(my_cos(2424)),16);
when x"979" => lut_sig <= to_unsigned(integer(my_cos(2425)),16);
when x"97a" => lut_sig <= to_unsigned(integer(my_cos(2426)),16);
when x"97b" => lut_sig <= to_unsigned(integer(my_cos(2427)),16);
when x"97c" => lut_sig <= to_unsigned(integer(my_cos(2428)),16);
when x"97d" => lut_sig <= to_unsigned(integer(my_cos(2429)),16);
when x"97e" => lut_sig <= to_unsigned(integer(my_cos(2430)),16);
when x"97f" => lut_sig <= to_unsigned(integer(my_cos(2431)),16);
when x"980" => lut_sig <= to_unsigned(integer(my_cos(2432)),16);
when x"981" => lut_sig <= to_unsigned(integer(my_cos(2433)),16);
when x"982" => lut_sig <= to_unsigned(integer(my_cos(2434)),16);
when x"983" => lut_sig <= to_unsigned(integer(my_cos(2435)),16);
when x"984" => lut_sig <= to_unsigned(integer(my_cos(2436)),16);
when x"985" => lut_sig <= to_unsigned(integer(my_cos(2437)),16);
when x"986" => lut_sig <= to_unsigned(integer(my_cos(2438)),16);
when x"987" => lut_sig <= to_unsigned(integer(my_cos(2439)),16);
when x"988" => lut_sig <= to_unsigned(integer(my_cos(2440)),16);
when x"989" => lut_sig <= to_unsigned(integer(my_cos(2441)),16);
when x"98a" => lut_sig <= to_unsigned(integer(my_cos(2442)),16);
when x"98b" => lut_sig <= to_unsigned(integer(my_cos(2443)),16);
when x"98c" => lut_sig <= to_unsigned(integer(my_cos(2444)),16);
when x"98d" => lut_sig <= to_unsigned(integer(my_cos(2445)),16);
when x"98e" => lut_sig <= to_unsigned(integer(my_cos(2446)),16);
when x"98f" => lut_sig <= to_unsigned(integer(my_cos(2447)),16);
when x"990" => lut_sig <= to_unsigned(integer(my_cos(2448)),16);
when x"991" => lut_sig <= to_unsigned(integer(my_cos(2449)),16);
when x"992" => lut_sig <= to_unsigned(integer(my_cos(2450)),16);
when x"993" => lut_sig <= to_unsigned(integer(my_cos(2451)),16);
when x"994" => lut_sig <= to_unsigned(integer(my_cos(2452)),16);
when x"995" => lut_sig <= to_unsigned(integer(my_cos(2453)),16);
when x"996" => lut_sig <= to_unsigned(integer(my_cos(2454)),16);
when x"997" => lut_sig <= to_unsigned(integer(my_cos(2455)),16);
when x"998" => lut_sig <= to_unsigned(integer(my_cos(2456)),16);
when x"999" => lut_sig <= to_unsigned(integer(my_cos(2457)),16);
when x"99a" => lut_sig <= to_unsigned(integer(my_cos(2458)),16);
when x"99b" => lut_sig <= to_unsigned(integer(my_cos(2459)),16);
when x"99c" => lut_sig <= to_unsigned(integer(my_cos(2460)),16);
when x"99d" => lut_sig <= to_unsigned(integer(my_cos(2461)),16);
when x"99e" => lut_sig <= to_unsigned(integer(my_cos(2462)),16);
when x"99f" => lut_sig <= to_unsigned(integer(my_cos(2463)),16);
when x"9a0" => lut_sig <= to_unsigned(integer(my_cos(2464)),16);
when x"9a1" => lut_sig <= to_unsigned(integer(my_cos(2465)),16);
when x"9a2" => lut_sig <= to_unsigned(integer(my_cos(2466)),16);
when x"9a3" => lut_sig <= to_unsigned(integer(my_cos(2467)),16);
when x"9a4" => lut_sig <= to_unsigned(integer(my_cos(2468)),16);
when x"9a5" => lut_sig <= to_unsigned(integer(my_cos(2469)),16);
when x"9a6" => lut_sig <= to_unsigned(integer(my_cos(2470)),16);
when x"9a7" => lut_sig <= to_unsigned(integer(my_cos(2471)),16);
when x"9a8" => lut_sig <= to_unsigned(integer(my_cos(2472)),16);
when x"9a9" => lut_sig <= to_unsigned(integer(my_cos(2473)),16);
when x"9aa" => lut_sig <= to_unsigned(integer(my_cos(2474)),16);
when x"9ab" => lut_sig <= to_unsigned(integer(my_cos(2475)),16);
when x"9ac" => lut_sig <= to_unsigned(integer(my_cos(2476)),16);
when x"9ad" => lut_sig <= to_unsigned(integer(my_cos(2477)),16);
when x"9ae" => lut_sig <= to_unsigned(integer(my_cos(2478)),16);
when x"9af" => lut_sig <= to_unsigned(integer(my_cos(2479)),16);
when x"9b0" => lut_sig <= to_unsigned(integer(my_cos(2480)),16);
when x"9b1" => lut_sig <= to_unsigned(integer(my_cos(2481)),16);
when x"9b2" => lut_sig <= to_unsigned(integer(my_cos(2482)),16);
when x"9b3" => lut_sig <= to_unsigned(integer(my_cos(2483)),16);
when x"9b4" => lut_sig <= to_unsigned(integer(my_cos(2484)),16);
when x"9b5" => lut_sig <= to_unsigned(integer(my_cos(2485)),16);
when x"9b6" => lut_sig <= to_unsigned(integer(my_cos(2486)),16);
when x"9b7" => lut_sig <= to_unsigned(integer(my_cos(2487)),16);
when x"9b8" => lut_sig <= to_unsigned(integer(my_cos(2488)),16);
when x"9b9" => lut_sig <= to_unsigned(integer(my_cos(2489)),16);
when x"9ba" => lut_sig <= to_unsigned(integer(my_cos(2490)),16);
when x"9bb" => lut_sig <= to_unsigned(integer(my_cos(2491)),16);
when x"9bc" => lut_sig <= to_unsigned(integer(my_cos(2492)),16);
when x"9bd" => lut_sig <= to_unsigned(integer(my_cos(2493)),16);
when x"9be" => lut_sig <= to_unsigned(integer(my_cos(2494)),16);
when x"9bf" => lut_sig <= to_unsigned(integer(my_cos(2495)),16);
when x"9c0" => lut_sig <= to_unsigned(integer(my_cos(2496)),16);
when x"9c1" => lut_sig <= to_unsigned(integer(my_cos(2497)),16);
when x"9c2" => lut_sig <= to_unsigned(integer(my_cos(2498)),16);
when x"9c3" => lut_sig <= to_unsigned(integer(my_cos(2499)),16);
when x"9c4" => lut_sig <= to_unsigned(integer(my_cos(2500)),16);
when x"9c5" => lut_sig <= to_unsigned(integer(my_cos(2501)),16);
when x"9c6" => lut_sig <= to_unsigned(integer(my_cos(2502)),16);
when x"9c7" => lut_sig <= to_unsigned(integer(my_cos(2503)),16);
when x"9c8" => lut_sig <= to_unsigned(integer(my_cos(2504)),16);
when x"9c9" => lut_sig <= to_unsigned(integer(my_cos(2505)),16);
when x"9ca" => lut_sig <= to_unsigned(integer(my_cos(2506)),16);
when x"9cb" => lut_sig <= to_unsigned(integer(my_cos(2507)),16);
when x"9cc" => lut_sig <= to_unsigned(integer(my_cos(2508)),16);
when x"9cd" => lut_sig <= to_unsigned(integer(my_cos(2509)),16);
when x"9ce" => lut_sig <= to_unsigned(integer(my_cos(2510)),16);
when x"9cf" => lut_sig <= to_unsigned(integer(my_cos(2511)),16);
when x"9d0" => lut_sig <= to_unsigned(integer(my_cos(2512)),16);
when x"9d1" => lut_sig <= to_unsigned(integer(my_cos(2513)),16);
when x"9d2" => lut_sig <= to_unsigned(integer(my_cos(2514)),16);
when x"9d3" => lut_sig <= to_unsigned(integer(my_cos(2515)),16);
when x"9d4" => lut_sig <= to_unsigned(integer(my_cos(2516)),16);
when x"9d5" => lut_sig <= to_unsigned(integer(my_cos(2517)),16);
when x"9d6" => lut_sig <= to_unsigned(integer(my_cos(2518)),16);
when x"9d7" => lut_sig <= to_unsigned(integer(my_cos(2519)),16);
when x"9d8" => lut_sig <= to_unsigned(integer(my_cos(2520)),16);
when x"9d9" => lut_sig <= to_unsigned(integer(my_cos(2521)),16);
when x"9da" => lut_sig <= to_unsigned(integer(my_cos(2522)),16);
when x"9db" => lut_sig <= to_unsigned(integer(my_cos(2523)),16);
when x"9dc" => lut_sig <= to_unsigned(integer(my_cos(2524)),16);
when x"9dd" => lut_sig <= to_unsigned(integer(my_cos(2525)),16);
when x"9de" => lut_sig <= to_unsigned(integer(my_cos(2526)),16);
when x"9df" => lut_sig <= to_unsigned(integer(my_cos(2527)),16);
when x"9e0" => lut_sig <= to_unsigned(integer(my_cos(2528)),16);
when x"9e1" => lut_sig <= to_unsigned(integer(my_cos(2529)),16);
when x"9e2" => lut_sig <= to_unsigned(integer(my_cos(2530)),16);
when x"9e3" => lut_sig <= to_unsigned(integer(my_cos(2531)),16);
when x"9e4" => lut_sig <= to_unsigned(integer(my_cos(2532)),16);
when x"9e5" => lut_sig <= to_unsigned(integer(my_cos(2533)),16);
when x"9e6" => lut_sig <= to_unsigned(integer(my_cos(2534)),16);
when x"9e7" => lut_sig <= to_unsigned(integer(my_cos(2535)),16);
when x"9e8" => lut_sig <= to_unsigned(integer(my_cos(2536)),16);
when x"9e9" => lut_sig <= to_unsigned(integer(my_cos(2537)),16);
when x"9ea" => lut_sig <= to_unsigned(integer(my_cos(2538)),16);
when x"9eb" => lut_sig <= to_unsigned(integer(my_cos(2539)),16);
when x"9ec" => lut_sig <= to_unsigned(integer(my_cos(2540)),16);
when x"9ed" => lut_sig <= to_unsigned(integer(my_cos(2541)),16);
when x"9ee" => lut_sig <= to_unsigned(integer(my_cos(2542)),16);
when x"9ef" => lut_sig <= to_unsigned(integer(my_cos(2543)),16);
when x"9f0" => lut_sig <= to_unsigned(integer(my_cos(2544)),16);
when x"9f1" => lut_sig <= to_unsigned(integer(my_cos(2545)),16);
when x"9f2" => lut_sig <= to_unsigned(integer(my_cos(2546)),16);
when x"9f3" => lut_sig <= to_unsigned(integer(my_cos(2547)),16);
when x"9f4" => lut_sig <= to_unsigned(integer(my_cos(2548)),16);
when x"9f5" => lut_sig <= to_unsigned(integer(my_cos(2549)),16);
when x"9f6" => lut_sig <= to_unsigned(integer(my_cos(2550)),16);
when x"9f7" => lut_sig <= to_unsigned(integer(my_cos(2551)),16);
when x"9f8" => lut_sig <= to_unsigned(integer(my_cos(2552)),16);
when x"9f9" => lut_sig <= to_unsigned(integer(my_cos(2553)),16);
when x"9fa" => lut_sig <= to_unsigned(integer(my_cos(2554)),16);
when x"9fb" => lut_sig <= to_unsigned(integer(my_cos(2555)),16);
when x"9fc" => lut_sig <= to_unsigned(integer(my_cos(2556)),16);
when x"9fd" => lut_sig <= to_unsigned(integer(my_cos(2557)),16);
when x"9fe" => lut_sig <= to_unsigned(integer(my_cos(2558)),16);
when x"9ff" => lut_sig <= to_unsigned(integer(my_cos(2559)),16);
when x"a00" => lut_sig <= to_unsigned(integer(my_cos(2560)),16);
when x"a01" => lut_sig <= to_unsigned(integer(my_cos(2561)),16);
when x"a02" => lut_sig <= to_unsigned(integer(my_cos(2562)),16);
when x"a03" => lut_sig <= to_unsigned(integer(my_cos(2563)),16);
when x"a04" => lut_sig <= to_unsigned(integer(my_cos(2564)),16);
when x"a05" => lut_sig <= to_unsigned(integer(my_cos(2565)),16);
when x"a06" => lut_sig <= to_unsigned(integer(my_cos(2566)),16);
when x"a07" => lut_sig <= to_unsigned(integer(my_cos(2567)),16);
when x"a08" => lut_sig <= to_unsigned(integer(my_cos(2568)),16);
when x"a09" => lut_sig <= to_unsigned(integer(my_cos(2569)),16);
when x"a0a" => lut_sig <= to_unsigned(integer(my_cos(2570)),16);
when x"a0b" => lut_sig <= to_unsigned(integer(my_cos(2571)),16);
when x"a0c" => lut_sig <= to_unsigned(integer(my_cos(2572)),16);
when x"a0d" => lut_sig <= to_unsigned(integer(my_cos(2573)),16);
when x"a0e" => lut_sig <= to_unsigned(integer(my_cos(2574)),16);
when x"a0f" => lut_sig <= to_unsigned(integer(my_cos(2575)),16);
when x"a10" => lut_sig <= to_unsigned(integer(my_cos(2576)),16);
when x"a11" => lut_sig <= to_unsigned(integer(my_cos(2577)),16);
when x"a12" => lut_sig <= to_unsigned(integer(my_cos(2578)),16);
when x"a13" => lut_sig <= to_unsigned(integer(my_cos(2579)),16);
when x"a14" => lut_sig <= to_unsigned(integer(my_cos(2580)),16);
when x"a15" => lut_sig <= to_unsigned(integer(my_cos(2581)),16);
when x"a16" => lut_sig <= to_unsigned(integer(my_cos(2582)),16);
when x"a17" => lut_sig <= to_unsigned(integer(my_cos(2583)),16);
when x"a18" => lut_sig <= to_unsigned(integer(my_cos(2584)),16);
when x"a19" => lut_sig <= to_unsigned(integer(my_cos(2585)),16);
when x"a1a" => lut_sig <= to_unsigned(integer(my_cos(2586)),16);
when x"a1b" => lut_sig <= to_unsigned(integer(my_cos(2587)),16);
when x"a1c" => lut_sig <= to_unsigned(integer(my_cos(2588)),16);
when x"a1d" => lut_sig <= to_unsigned(integer(my_cos(2589)),16);
when x"a1e" => lut_sig <= to_unsigned(integer(my_cos(2590)),16);
when x"a1f" => lut_sig <= to_unsigned(integer(my_cos(2591)),16);
when x"a20" => lut_sig <= to_unsigned(integer(my_cos(2592)),16);
when x"a21" => lut_sig <= to_unsigned(integer(my_cos(2593)),16);
when x"a22" => lut_sig <= to_unsigned(integer(my_cos(2594)),16);
when x"a23" => lut_sig <= to_unsigned(integer(my_cos(2595)),16);
when x"a24" => lut_sig <= to_unsigned(integer(my_cos(2596)),16);
when x"a25" => lut_sig <= to_unsigned(integer(my_cos(2597)),16);
when x"a26" => lut_sig <= to_unsigned(integer(my_cos(2598)),16);
when x"a27" => lut_sig <= to_unsigned(integer(my_cos(2599)),16);
when x"a28" => lut_sig <= to_unsigned(integer(my_cos(2600)),16);
when x"a29" => lut_sig <= to_unsigned(integer(my_cos(2601)),16);
when x"a2a" => lut_sig <= to_unsigned(integer(my_cos(2602)),16);
when x"a2b" => lut_sig <= to_unsigned(integer(my_cos(2603)),16);
when x"a2c" => lut_sig <= to_unsigned(integer(my_cos(2604)),16);
when x"a2d" => lut_sig <= to_unsigned(integer(my_cos(2605)),16);
when x"a2e" => lut_sig <= to_unsigned(integer(my_cos(2606)),16);
when x"a2f" => lut_sig <= to_unsigned(integer(my_cos(2607)),16);
when x"a30" => lut_sig <= to_unsigned(integer(my_cos(2608)),16);
when x"a31" => lut_sig <= to_unsigned(integer(my_cos(2609)),16);
when x"a32" => lut_sig <= to_unsigned(integer(my_cos(2610)),16);
when x"a33" => lut_sig <= to_unsigned(integer(my_cos(2611)),16);
when x"a34" => lut_sig <= to_unsigned(integer(my_cos(2612)),16);
when x"a35" => lut_sig <= to_unsigned(integer(my_cos(2613)),16);
when x"a36" => lut_sig <= to_unsigned(integer(my_cos(2614)),16);
when x"a37" => lut_sig <= to_unsigned(integer(my_cos(2615)),16);
when x"a38" => lut_sig <= to_unsigned(integer(my_cos(2616)),16);
when x"a39" => lut_sig <= to_unsigned(integer(my_cos(2617)),16);
when x"a3a" => lut_sig <= to_unsigned(integer(my_cos(2618)),16);
when x"a3b" => lut_sig <= to_unsigned(integer(my_cos(2619)),16);
when x"a3c" => lut_sig <= to_unsigned(integer(my_cos(2620)),16);
when x"a3d" => lut_sig <= to_unsigned(integer(my_cos(2621)),16);
when x"a3e" => lut_sig <= to_unsigned(integer(my_cos(2622)),16);
when x"a3f" => lut_sig <= to_unsigned(integer(my_cos(2623)),16);
when x"a40" => lut_sig <= to_unsigned(integer(my_cos(2624)),16);
when x"a41" => lut_sig <= to_unsigned(integer(my_cos(2625)),16);
when x"a42" => lut_sig <= to_unsigned(integer(my_cos(2626)),16);
when x"a43" => lut_sig <= to_unsigned(integer(my_cos(2627)),16);
when x"a44" => lut_sig <= to_unsigned(integer(my_cos(2628)),16);
when x"a45" => lut_sig <= to_unsigned(integer(my_cos(2629)),16);
when x"a46" => lut_sig <= to_unsigned(integer(my_cos(2630)),16);
when x"a47" => lut_sig <= to_unsigned(integer(my_cos(2631)),16);
when x"a48" => lut_sig <= to_unsigned(integer(my_cos(2632)),16);
when x"a49" => lut_sig <= to_unsigned(integer(my_cos(2633)),16);
when x"a4a" => lut_sig <= to_unsigned(integer(my_cos(2634)),16);
when x"a4b" => lut_sig <= to_unsigned(integer(my_cos(2635)),16);
when x"a4c" => lut_sig <= to_unsigned(integer(my_cos(2636)),16);
when x"a4d" => lut_sig <= to_unsigned(integer(my_cos(2637)),16);
when x"a4e" => lut_sig <= to_unsigned(integer(my_cos(2638)),16);
when x"a4f" => lut_sig <= to_unsigned(integer(my_cos(2639)),16);
when x"a50" => lut_sig <= to_unsigned(integer(my_cos(2640)),16);
when x"a51" => lut_sig <= to_unsigned(integer(my_cos(2641)),16);
when x"a52" => lut_sig <= to_unsigned(integer(my_cos(2642)),16);
when x"a53" => lut_sig <= to_unsigned(integer(my_cos(2643)),16);
when x"a54" => lut_sig <= to_unsigned(integer(my_cos(2644)),16);
when x"a55" => lut_sig <= to_unsigned(integer(my_cos(2645)),16);
when x"a56" => lut_sig <= to_unsigned(integer(my_cos(2646)),16);
when x"a57" => lut_sig <= to_unsigned(integer(my_cos(2647)),16);
when x"a58" => lut_sig <= to_unsigned(integer(my_cos(2648)),16);
when x"a59" => lut_sig <= to_unsigned(integer(my_cos(2649)),16);
when x"a5a" => lut_sig <= to_unsigned(integer(my_cos(2650)),16);
when x"a5b" => lut_sig <= to_unsigned(integer(my_cos(2651)),16);
when x"a5c" => lut_sig <= to_unsigned(integer(my_cos(2652)),16);
when x"a5d" => lut_sig <= to_unsigned(integer(my_cos(2653)),16);
when x"a5e" => lut_sig <= to_unsigned(integer(my_cos(2654)),16);
when x"a5f" => lut_sig <= to_unsigned(integer(my_cos(2655)),16);
when x"a60" => lut_sig <= to_unsigned(integer(my_cos(2656)),16);
when x"a61" => lut_sig <= to_unsigned(integer(my_cos(2657)),16);
when x"a62" => lut_sig <= to_unsigned(integer(my_cos(2658)),16);
when x"a63" => lut_sig <= to_unsigned(integer(my_cos(2659)),16);
when x"a64" => lut_sig <= to_unsigned(integer(my_cos(2660)),16);
when x"a65" => lut_sig <= to_unsigned(integer(my_cos(2661)),16);
when x"a66" => lut_sig <= to_unsigned(integer(my_cos(2662)),16);
when x"a67" => lut_sig <= to_unsigned(integer(my_cos(2663)),16);
when x"a68" => lut_sig <= to_unsigned(integer(my_cos(2664)),16);
when x"a69" => lut_sig <= to_unsigned(integer(my_cos(2665)),16);
when x"a6a" => lut_sig <= to_unsigned(integer(my_cos(2666)),16);
when x"a6b" => lut_sig <= to_unsigned(integer(my_cos(2667)),16);
when x"a6c" => lut_sig <= to_unsigned(integer(my_cos(2668)),16);
when x"a6d" => lut_sig <= to_unsigned(integer(my_cos(2669)),16);
when x"a6e" => lut_sig <= to_unsigned(integer(my_cos(2670)),16);
when x"a6f" => lut_sig <= to_unsigned(integer(my_cos(2671)),16);
when x"a70" => lut_sig <= to_unsigned(integer(my_cos(2672)),16);
when x"a71" => lut_sig <= to_unsigned(integer(my_cos(2673)),16);
when x"a72" => lut_sig <= to_unsigned(integer(my_cos(2674)),16);
when x"a73" => lut_sig <= to_unsigned(integer(my_cos(2675)),16);
when x"a74" => lut_sig <= to_unsigned(integer(my_cos(2676)),16);
when x"a75" => lut_sig <= to_unsigned(integer(my_cos(2677)),16);
when x"a76" => lut_sig <= to_unsigned(integer(my_cos(2678)),16);
when x"a77" => lut_sig <= to_unsigned(integer(my_cos(2679)),16);
when x"a78" => lut_sig <= to_unsigned(integer(my_cos(2680)),16);
when x"a79" => lut_sig <= to_unsigned(integer(my_cos(2681)),16);
when x"a7a" => lut_sig <= to_unsigned(integer(my_cos(2682)),16);
when x"a7b" => lut_sig <= to_unsigned(integer(my_cos(2683)),16);
when x"a7c" => lut_sig <= to_unsigned(integer(my_cos(2684)),16);
when x"a7d" => lut_sig <= to_unsigned(integer(my_cos(2685)),16);
when x"a7e" => lut_sig <= to_unsigned(integer(my_cos(2686)),16);
when x"a7f" => lut_sig <= to_unsigned(integer(my_cos(2687)),16);
when x"a80" => lut_sig <= to_unsigned(integer(my_cos(2688)),16);
when x"a81" => lut_sig <= to_unsigned(integer(my_cos(2689)),16);
when x"a82" => lut_sig <= to_unsigned(integer(my_cos(2690)),16);
when x"a83" => lut_sig <= to_unsigned(integer(my_cos(2691)),16);
when x"a84" => lut_sig <= to_unsigned(integer(my_cos(2692)),16);
when x"a85" => lut_sig <= to_unsigned(integer(my_cos(2693)),16);
when x"a86" => lut_sig <= to_unsigned(integer(my_cos(2694)),16);
when x"a87" => lut_sig <= to_unsigned(integer(my_cos(2695)),16);
when x"a88" => lut_sig <= to_unsigned(integer(my_cos(2696)),16);
when x"a89" => lut_sig <= to_unsigned(integer(my_cos(2697)),16);
when x"a8a" => lut_sig <= to_unsigned(integer(my_cos(2698)),16);
when x"a8b" => lut_sig <= to_unsigned(integer(my_cos(2699)),16);
when x"a8c" => lut_sig <= to_unsigned(integer(my_cos(2700)),16);
when x"a8d" => lut_sig <= to_unsigned(integer(my_cos(2701)),16);
when x"a8e" => lut_sig <= to_unsigned(integer(my_cos(2702)),16);
when x"a8f" => lut_sig <= to_unsigned(integer(my_cos(2703)),16);
when x"a90" => lut_sig <= to_unsigned(integer(my_cos(2704)),16);
when x"a91" => lut_sig <= to_unsigned(integer(my_cos(2705)),16);
when x"a92" => lut_sig <= to_unsigned(integer(my_cos(2706)),16);
when x"a93" => lut_sig <= to_unsigned(integer(my_cos(2707)),16);
when x"a94" => lut_sig <= to_unsigned(integer(my_cos(2708)),16);
when x"a95" => lut_sig <= to_unsigned(integer(my_cos(2709)),16);
when x"a96" => lut_sig <= to_unsigned(integer(my_cos(2710)),16);
when x"a97" => lut_sig <= to_unsigned(integer(my_cos(2711)),16);
when x"a98" => lut_sig <= to_unsigned(integer(my_cos(2712)),16);
when x"a99" => lut_sig <= to_unsigned(integer(my_cos(2713)),16);
when x"a9a" => lut_sig <= to_unsigned(integer(my_cos(2714)),16);
when x"a9b" => lut_sig <= to_unsigned(integer(my_cos(2715)),16);
when x"a9c" => lut_sig <= to_unsigned(integer(my_cos(2716)),16);
when x"a9d" => lut_sig <= to_unsigned(integer(my_cos(2717)),16);
when x"a9e" => lut_sig <= to_unsigned(integer(my_cos(2718)),16);
when x"a9f" => lut_sig <= to_unsigned(integer(my_cos(2719)),16);
when x"aa0" => lut_sig <= to_unsigned(integer(my_cos(2720)),16);
when x"aa1" => lut_sig <= to_unsigned(integer(my_cos(2721)),16);
when x"aa2" => lut_sig <= to_unsigned(integer(my_cos(2722)),16);
when x"aa3" => lut_sig <= to_unsigned(integer(my_cos(2723)),16);
when x"aa4" => lut_sig <= to_unsigned(integer(my_cos(2724)),16);
when x"aa5" => lut_sig <= to_unsigned(integer(my_cos(2725)),16);
when x"aa6" => lut_sig <= to_unsigned(integer(my_cos(2726)),16);
when x"aa7" => lut_sig <= to_unsigned(integer(my_cos(2727)),16);
when x"aa8" => lut_sig <= to_unsigned(integer(my_cos(2728)),16);
when x"aa9" => lut_sig <= to_unsigned(integer(my_cos(2729)),16);
when x"aaa" => lut_sig <= to_unsigned(integer(my_cos(2730)),16);
when x"aab" => lut_sig <= to_unsigned(integer(my_cos(2731)),16);
when x"aac" => lut_sig <= to_unsigned(integer(my_cos(2732)),16);
when x"aad" => lut_sig <= to_unsigned(integer(my_cos(2733)),16);
when x"aae" => lut_sig <= to_unsigned(integer(my_cos(2734)),16);
when x"aaf" => lut_sig <= to_unsigned(integer(my_cos(2735)),16);
when x"ab0" => lut_sig <= to_unsigned(integer(my_cos(2736)),16);
when x"ab1" => lut_sig <= to_unsigned(integer(my_cos(2737)),16);
when x"ab2" => lut_sig <= to_unsigned(integer(my_cos(2738)),16);
when x"ab3" => lut_sig <= to_unsigned(integer(my_cos(2739)),16);
when x"ab4" => lut_sig <= to_unsigned(integer(my_cos(2740)),16);
when x"ab5" => lut_sig <= to_unsigned(integer(my_cos(2741)),16);
when x"ab6" => lut_sig <= to_unsigned(integer(my_cos(2742)),16);
when x"ab7" => lut_sig <= to_unsigned(integer(my_cos(2743)),16);
when x"ab8" => lut_sig <= to_unsigned(integer(my_cos(2744)),16);
when x"ab9" => lut_sig <= to_unsigned(integer(my_cos(2745)),16);
when x"aba" => lut_sig <= to_unsigned(integer(my_cos(2746)),16);
when x"abb" => lut_sig <= to_unsigned(integer(my_cos(2747)),16);
when x"abc" => lut_sig <= to_unsigned(integer(my_cos(2748)),16);
when x"abd" => lut_sig <= to_unsigned(integer(my_cos(2749)),16);
when x"abe" => lut_sig <= to_unsigned(integer(my_cos(2750)),16);
when x"abf" => lut_sig <= to_unsigned(integer(my_cos(2751)),16);
when x"ac0" => lut_sig <= to_unsigned(integer(my_cos(2752)),16);
when x"ac1" => lut_sig <= to_unsigned(integer(my_cos(2753)),16);
when x"ac2" => lut_sig <= to_unsigned(integer(my_cos(2754)),16);
when x"ac3" => lut_sig <= to_unsigned(integer(my_cos(2755)),16);
when x"ac4" => lut_sig <= to_unsigned(integer(my_cos(2756)),16);
when x"ac5" => lut_sig <= to_unsigned(integer(my_cos(2757)),16);
when x"ac6" => lut_sig <= to_unsigned(integer(my_cos(2758)),16);
when x"ac7" => lut_sig <= to_unsigned(integer(my_cos(2759)),16);
when x"ac8" => lut_sig <= to_unsigned(integer(my_cos(2760)),16);
when x"ac9" => lut_sig <= to_unsigned(integer(my_cos(2761)),16);
when x"aca" => lut_sig <= to_unsigned(integer(my_cos(2762)),16);
when x"acb" => lut_sig <= to_unsigned(integer(my_cos(2763)),16);
when x"acc" => lut_sig <= to_unsigned(integer(my_cos(2764)),16);
when x"acd" => lut_sig <= to_unsigned(integer(my_cos(2765)),16);
when x"ace" => lut_sig <= to_unsigned(integer(my_cos(2766)),16);
when x"acf" => lut_sig <= to_unsigned(integer(my_cos(2767)),16);
when x"ad0" => lut_sig <= to_unsigned(integer(my_cos(2768)),16);
when x"ad1" => lut_sig <= to_unsigned(integer(my_cos(2769)),16);
when x"ad2" => lut_sig <= to_unsigned(integer(my_cos(2770)),16);
when x"ad3" => lut_sig <= to_unsigned(integer(my_cos(2771)),16);
when x"ad4" => lut_sig <= to_unsigned(integer(my_cos(2772)),16);
when x"ad5" => lut_sig <= to_unsigned(integer(my_cos(2773)),16);
when x"ad6" => lut_sig <= to_unsigned(integer(my_cos(2774)),16);
when x"ad7" => lut_sig <= to_unsigned(integer(my_cos(2775)),16);
when x"ad8" => lut_sig <= to_unsigned(integer(my_cos(2776)),16);
when x"ad9" => lut_sig <= to_unsigned(integer(my_cos(2777)),16);
when x"ada" => lut_sig <= to_unsigned(integer(my_cos(2778)),16);
when x"adb" => lut_sig <= to_unsigned(integer(my_cos(2779)),16);
when x"adc" => lut_sig <= to_unsigned(integer(my_cos(2780)),16);
when x"add" => lut_sig <= to_unsigned(integer(my_cos(2781)),16);
when x"ade" => lut_sig <= to_unsigned(integer(my_cos(2782)),16);
when x"adf" => lut_sig <= to_unsigned(integer(my_cos(2783)),16);
when x"ae0" => lut_sig <= to_unsigned(integer(my_cos(2784)),16);
when x"ae1" => lut_sig <= to_unsigned(integer(my_cos(2785)),16);
when x"ae2" => lut_sig <= to_unsigned(integer(my_cos(2786)),16);
when x"ae3" => lut_sig <= to_unsigned(integer(my_cos(2787)),16);
when x"ae4" => lut_sig <= to_unsigned(integer(my_cos(2788)),16);
when x"ae5" => lut_sig <= to_unsigned(integer(my_cos(2789)),16);
when x"ae6" => lut_sig <= to_unsigned(integer(my_cos(2790)),16);
when x"ae7" => lut_sig <= to_unsigned(integer(my_cos(2791)),16);
when x"ae8" => lut_sig <= to_unsigned(integer(my_cos(2792)),16);
when x"ae9" => lut_sig <= to_unsigned(integer(my_cos(2793)),16);
when x"aea" => lut_sig <= to_unsigned(integer(my_cos(2794)),16);
when x"aeb" => lut_sig <= to_unsigned(integer(my_cos(2795)),16);
when x"aec" => lut_sig <= to_unsigned(integer(my_cos(2796)),16);
when x"aed" => lut_sig <= to_unsigned(integer(my_cos(2797)),16);
when x"aee" => lut_sig <= to_unsigned(integer(my_cos(2798)),16);
when x"aef" => lut_sig <= to_unsigned(integer(my_cos(2799)),16);
when x"af0" => lut_sig <= to_unsigned(integer(my_cos(2800)),16);
when x"af1" => lut_sig <= to_unsigned(integer(my_cos(2801)),16);
when x"af2" => lut_sig <= to_unsigned(integer(my_cos(2802)),16);
when x"af3" => lut_sig <= to_unsigned(integer(my_cos(2803)),16);
when x"af4" => lut_sig <= to_unsigned(integer(my_cos(2804)),16);
when x"af5" => lut_sig <= to_unsigned(integer(my_cos(2805)),16);
when x"af6" => lut_sig <= to_unsigned(integer(my_cos(2806)),16);
when x"af7" => lut_sig <= to_unsigned(integer(my_cos(2807)),16);
when x"af8" => lut_sig <= to_unsigned(integer(my_cos(2808)),16);
when x"af9" => lut_sig <= to_unsigned(integer(my_cos(2809)),16);
when x"afa" => lut_sig <= to_unsigned(integer(my_cos(2810)),16);
when x"afb" => lut_sig <= to_unsigned(integer(my_cos(2811)),16);
when x"afc" => lut_sig <= to_unsigned(integer(my_cos(2812)),16);
when x"afd" => lut_sig <= to_unsigned(integer(my_cos(2813)),16);
when x"afe" => lut_sig <= to_unsigned(integer(my_cos(2814)),16);
when x"aff" => lut_sig <= to_unsigned(integer(my_cos(2815)),16);
when x"b00" => lut_sig <= to_unsigned(integer(my_cos(2816)),16);
when x"b01" => lut_sig <= to_unsigned(integer(my_cos(2817)),16);
when x"b02" => lut_sig <= to_unsigned(integer(my_cos(2818)),16);
when x"b03" => lut_sig <= to_unsigned(integer(my_cos(2819)),16);
when x"b04" => lut_sig <= to_unsigned(integer(my_cos(2820)),16);
when x"b05" => lut_sig <= to_unsigned(integer(my_cos(2821)),16);
when x"b06" => lut_sig <= to_unsigned(integer(my_cos(2822)),16);
when x"b07" => lut_sig <= to_unsigned(integer(my_cos(2823)),16);
when x"b08" => lut_sig <= to_unsigned(integer(my_cos(2824)),16);
when x"b09" => lut_sig <= to_unsigned(integer(my_cos(2825)),16);
when x"b0a" => lut_sig <= to_unsigned(integer(my_cos(2826)),16);
when x"b0b" => lut_sig <= to_unsigned(integer(my_cos(2827)),16);
when x"b0c" => lut_sig <= to_unsigned(integer(my_cos(2828)),16);
when x"b0d" => lut_sig <= to_unsigned(integer(my_cos(2829)),16);
when x"b0e" => lut_sig <= to_unsigned(integer(my_cos(2830)),16);
when x"b0f" => lut_sig <= to_unsigned(integer(my_cos(2831)),16);
when x"b10" => lut_sig <= to_unsigned(integer(my_cos(2832)),16);
when x"b11" => lut_sig <= to_unsigned(integer(my_cos(2833)),16);
when x"b12" => lut_sig <= to_unsigned(integer(my_cos(2834)),16);
when x"b13" => lut_sig <= to_unsigned(integer(my_cos(2835)),16);
when x"b14" => lut_sig <= to_unsigned(integer(my_cos(2836)),16);
when x"b15" => lut_sig <= to_unsigned(integer(my_cos(2837)),16);
when x"b16" => lut_sig <= to_unsigned(integer(my_cos(2838)),16);
when x"b17" => lut_sig <= to_unsigned(integer(my_cos(2839)),16);
when x"b18" => lut_sig <= to_unsigned(integer(my_cos(2840)),16);
when x"b19" => lut_sig <= to_unsigned(integer(my_cos(2841)),16);
when x"b1a" => lut_sig <= to_unsigned(integer(my_cos(2842)),16);
when x"b1b" => lut_sig <= to_unsigned(integer(my_cos(2843)),16);
when x"b1c" => lut_sig <= to_unsigned(integer(my_cos(2844)),16);
when x"b1d" => lut_sig <= to_unsigned(integer(my_cos(2845)),16);
when x"b1e" => lut_sig <= to_unsigned(integer(my_cos(2846)),16);
when x"b1f" => lut_sig <= to_unsigned(integer(my_cos(2847)),16);
when x"b20" => lut_sig <= to_unsigned(integer(my_cos(2848)),16);
when x"b21" => lut_sig <= to_unsigned(integer(my_cos(2849)),16);
when x"b22" => lut_sig <= to_unsigned(integer(my_cos(2850)),16);
when x"b23" => lut_sig <= to_unsigned(integer(my_cos(2851)),16);
when x"b24" => lut_sig <= to_unsigned(integer(my_cos(2852)),16);
when x"b25" => lut_sig <= to_unsigned(integer(my_cos(2853)),16);
when x"b26" => lut_sig <= to_unsigned(integer(my_cos(2854)),16);
when x"b27" => lut_sig <= to_unsigned(integer(my_cos(2855)),16);
when x"b28" => lut_sig <= to_unsigned(integer(my_cos(2856)),16);
when x"b29" => lut_sig <= to_unsigned(integer(my_cos(2857)),16);
when x"b2a" => lut_sig <= to_unsigned(integer(my_cos(2858)),16);
when x"b2b" => lut_sig <= to_unsigned(integer(my_cos(2859)),16);
when x"b2c" => lut_sig <= to_unsigned(integer(my_cos(2860)),16);
when x"b2d" => lut_sig <= to_unsigned(integer(my_cos(2861)),16);
when x"b2e" => lut_sig <= to_unsigned(integer(my_cos(2862)),16);
when x"b2f" => lut_sig <= to_unsigned(integer(my_cos(2863)),16);
when x"b30" => lut_sig <= to_unsigned(integer(my_cos(2864)),16);
when x"b31" => lut_sig <= to_unsigned(integer(my_cos(2865)),16);
when x"b32" => lut_sig <= to_unsigned(integer(my_cos(2866)),16);
when x"b33" => lut_sig <= to_unsigned(integer(my_cos(2867)),16);
when x"b34" => lut_sig <= to_unsigned(integer(my_cos(2868)),16);
when x"b35" => lut_sig <= to_unsigned(integer(my_cos(2869)),16);
when x"b36" => lut_sig <= to_unsigned(integer(my_cos(2870)),16);
when x"b37" => lut_sig <= to_unsigned(integer(my_cos(2871)),16);
when x"b38" => lut_sig <= to_unsigned(integer(my_cos(2872)),16);
when x"b39" => lut_sig <= to_unsigned(integer(my_cos(2873)),16);
when x"b3a" => lut_sig <= to_unsigned(integer(my_cos(2874)),16);
when x"b3b" => lut_sig <= to_unsigned(integer(my_cos(2875)),16);
when x"b3c" => lut_sig <= to_unsigned(integer(my_cos(2876)),16);
when x"b3d" => lut_sig <= to_unsigned(integer(my_cos(2877)),16);
when x"b3e" => lut_sig <= to_unsigned(integer(my_cos(2878)),16);
when x"b3f" => lut_sig <= to_unsigned(integer(my_cos(2879)),16);
when x"b40" => lut_sig <= to_unsigned(integer(my_cos(2880)),16);
when x"b41" => lut_sig <= to_unsigned(integer(my_cos(2881)),16);
when x"b42" => lut_sig <= to_unsigned(integer(my_cos(2882)),16);
when x"b43" => lut_sig <= to_unsigned(integer(my_cos(2883)),16);
when x"b44" => lut_sig <= to_unsigned(integer(my_cos(2884)),16);
when x"b45" => lut_sig <= to_unsigned(integer(my_cos(2885)),16);
when x"b46" => lut_sig <= to_unsigned(integer(my_cos(2886)),16);
when x"b47" => lut_sig <= to_unsigned(integer(my_cos(2887)),16);
when x"b48" => lut_sig <= to_unsigned(integer(my_cos(2888)),16);
when x"b49" => lut_sig <= to_unsigned(integer(my_cos(2889)),16);
when x"b4a" => lut_sig <= to_unsigned(integer(my_cos(2890)),16);
when x"b4b" => lut_sig <= to_unsigned(integer(my_cos(2891)),16);
when x"b4c" => lut_sig <= to_unsigned(integer(my_cos(2892)),16);
when x"b4d" => lut_sig <= to_unsigned(integer(my_cos(2893)),16);
when x"b4e" => lut_sig <= to_unsigned(integer(my_cos(2894)),16);
when x"b4f" => lut_sig <= to_unsigned(integer(my_cos(2895)),16);
when x"b50" => lut_sig <= to_unsigned(integer(my_cos(2896)),16);
when x"b51" => lut_sig <= to_unsigned(integer(my_cos(2897)),16);
when x"b52" => lut_sig <= to_unsigned(integer(my_cos(2898)),16);
when x"b53" => lut_sig <= to_unsigned(integer(my_cos(2899)),16);
when x"b54" => lut_sig <= to_unsigned(integer(my_cos(2900)),16);
when x"b55" => lut_sig <= to_unsigned(integer(my_cos(2901)),16);
when x"b56" => lut_sig <= to_unsigned(integer(my_cos(2902)),16);
when x"b57" => lut_sig <= to_unsigned(integer(my_cos(2903)),16);
when x"b58" => lut_sig <= to_unsigned(integer(my_cos(2904)),16);
when x"b59" => lut_sig <= to_unsigned(integer(my_cos(2905)),16);
when x"b5a" => lut_sig <= to_unsigned(integer(my_cos(2906)),16);
when x"b5b" => lut_sig <= to_unsigned(integer(my_cos(2907)),16);
when x"b5c" => lut_sig <= to_unsigned(integer(my_cos(2908)),16);
when x"b5d" => lut_sig <= to_unsigned(integer(my_cos(2909)),16);
when x"b5e" => lut_sig <= to_unsigned(integer(my_cos(2910)),16);
when x"b5f" => lut_sig <= to_unsigned(integer(my_cos(2911)),16);
when x"b60" => lut_sig <= to_unsigned(integer(my_cos(2912)),16);
when x"b61" => lut_sig <= to_unsigned(integer(my_cos(2913)),16);
when x"b62" => lut_sig <= to_unsigned(integer(my_cos(2914)),16);
when x"b63" => lut_sig <= to_unsigned(integer(my_cos(2915)),16);
when x"b64" => lut_sig <= to_unsigned(integer(my_cos(2916)),16);
when x"b65" => lut_sig <= to_unsigned(integer(my_cos(2917)),16);
when x"b66" => lut_sig <= to_unsigned(integer(my_cos(2918)),16);
when x"b67" => lut_sig <= to_unsigned(integer(my_cos(2919)),16);
when x"b68" => lut_sig <= to_unsigned(integer(my_cos(2920)),16);
when x"b69" => lut_sig <= to_unsigned(integer(my_cos(2921)),16);
when x"b6a" => lut_sig <= to_unsigned(integer(my_cos(2922)),16);
when x"b6b" => lut_sig <= to_unsigned(integer(my_cos(2923)),16);
when x"b6c" => lut_sig <= to_unsigned(integer(my_cos(2924)),16);
when x"b6d" => lut_sig <= to_unsigned(integer(my_cos(2925)),16);
when x"b6e" => lut_sig <= to_unsigned(integer(my_cos(2926)),16);
when x"b6f" => lut_sig <= to_unsigned(integer(my_cos(2927)),16);
when x"b70" => lut_sig <= to_unsigned(integer(my_cos(2928)),16);
when x"b71" => lut_sig <= to_unsigned(integer(my_cos(2929)),16);
when x"b72" => lut_sig <= to_unsigned(integer(my_cos(2930)),16);
when x"b73" => lut_sig <= to_unsigned(integer(my_cos(2931)),16);
when x"b74" => lut_sig <= to_unsigned(integer(my_cos(2932)),16);
when x"b75" => lut_sig <= to_unsigned(integer(my_cos(2933)),16);
when x"b76" => lut_sig <= to_unsigned(integer(my_cos(2934)),16);
when x"b77" => lut_sig <= to_unsigned(integer(my_cos(2935)),16);
when x"b78" => lut_sig <= to_unsigned(integer(my_cos(2936)),16);
when x"b79" => lut_sig <= to_unsigned(integer(my_cos(2937)),16);
when x"b7a" => lut_sig <= to_unsigned(integer(my_cos(2938)),16);
when x"b7b" => lut_sig <= to_unsigned(integer(my_cos(2939)),16);
when x"b7c" => lut_sig <= to_unsigned(integer(my_cos(2940)),16);
when x"b7d" => lut_sig <= to_unsigned(integer(my_cos(2941)),16);
when x"b7e" => lut_sig <= to_unsigned(integer(my_cos(2942)),16);
when x"b7f" => lut_sig <= to_unsigned(integer(my_cos(2943)),16);
when x"b80" => lut_sig <= to_unsigned(integer(my_cos(2944)),16);
when x"b81" => lut_sig <= to_unsigned(integer(my_cos(2945)),16);
when x"b82" => lut_sig <= to_unsigned(integer(my_cos(2946)),16);
when x"b83" => lut_sig <= to_unsigned(integer(my_cos(2947)),16);
when x"b84" => lut_sig <= to_unsigned(integer(my_cos(2948)),16);
when x"b85" => lut_sig <= to_unsigned(integer(my_cos(2949)),16);
when x"b86" => lut_sig <= to_unsigned(integer(my_cos(2950)),16);
when x"b87" => lut_sig <= to_unsigned(integer(my_cos(2951)),16);
when x"b88" => lut_sig <= to_unsigned(integer(my_cos(2952)),16);
when x"b89" => lut_sig <= to_unsigned(integer(my_cos(2953)),16);
when x"b8a" => lut_sig <= to_unsigned(integer(my_cos(2954)),16);
when x"b8b" => lut_sig <= to_unsigned(integer(my_cos(2955)),16);
when x"b8c" => lut_sig <= to_unsigned(integer(my_cos(2956)),16);
when x"b8d" => lut_sig <= to_unsigned(integer(my_cos(2957)),16);
when x"b8e" => lut_sig <= to_unsigned(integer(my_cos(2958)),16);
when x"b8f" => lut_sig <= to_unsigned(integer(my_cos(2959)),16);
when x"b90" => lut_sig <= to_unsigned(integer(my_cos(2960)),16);
when x"b91" => lut_sig <= to_unsigned(integer(my_cos(2961)),16);
when x"b92" => lut_sig <= to_unsigned(integer(my_cos(2962)),16);
when x"b93" => lut_sig <= to_unsigned(integer(my_cos(2963)),16);
when x"b94" => lut_sig <= to_unsigned(integer(my_cos(2964)),16);
when x"b95" => lut_sig <= to_unsigned(integer(my_cos(2965)),16);
when x"b96" => lut_sig <= to_unsigned(integer(my_cos(2966)),16);
when x"b97" => lut_sig <= to_unsigned(integer(my_cos(2967)),16);
when x"b98" => lut_sig <= to_unsigned(integer(my_cos(2968)),16);
when x"b99" => lut_sig <= to_unsigned(integer(my_cos(2969)),16);
when x"b9a" => lut_sig <= to_unsigned(integer(my_cos(2970)),16);
when x"b9b" => lut_sig <= to_unsigned(integer(my_cos(2971)),16);
when x"b9c" => lut_sig <= to_unsigned(integer(my_cos(2972)),16);
when x"b9d" => lut_sig <= to_unsigned(integer(my_cos(2973)),16);
when x"b9e" => lut_sig <= to_unsigned(integer(my_cos(2974)),16);
when x"b9f" => lut_sig <= to_unsigned(integer(my_cos(2975)),16);
when x"ba0" => lut_sig <= to_unsigned(integer(my_cos(2976)),16);
when x"ba1" => lut_sig <= to_unsigned(integer(my_cos(2977)),16);
when x"ba2" => lut_sig <= to_unsigned(integer(my_cos(2978)),16);
when x"ba3" => lut_sig <= to_unsigned(integer(my_cos(2979)),16);
when x"ba4" => lut_sig <= to_unsigned(integer(my_cos(2980)),16);
when x"ba5" => lut_sig <= to_unsigned(integer(my_cos(2981)),16);
when x"ba6" => lut_sig <= to_unsigned(integer(my_cos(2982)),16);
when x"ba7" => lut_sig <= to_unsigned(integer(my_cos(2983)),16);
when x"ba8" => lut_sig <= to_unsigned(integer(my_cos(2984)),16);
when x"ba9" => lut_sig <= to_unsigned(integer(my_cos(2985)),16);
when x"baa" => lut_sig <= to_unsigned(integer(my_cos(2986)),16);
when x"bab" => lut_sig <= to_unsigned(integer(my_cos(2987)),16);
when x"bac" => lut_sig <= to_unsigned(integer(my_cos(2988)),16);
when x"bad" => lut_sig <= to_unsigned(integer(my_cos(2989)),16);
when x"bae" => lut_sig <= to_unsigned(integer(my_cos(2990)),16);
when x"baf" => lut_sig <= to_unsigned(integer(my_cos(2991)),16);
when x"bb0" => lut_sig <= to_unsigned(integer(my_cos(2992)),16);
when x"bb1" => lut_sig <= to_unsigned(integer(my_cos(2993)),16);
when x"bb2" => lut_sig <= to_unsigned(integer(my_cos(2994)),16);
when x"bb3" => lut_sig <= to_unsigned(integer(my_cos(2995)),16);
when x"bb4" => lut_sig <= to_unsigned(integer(my_cos(2996)),16);
when x"bb5" => lut_sig <= to_unsigned(integer(my_cos(2997)),16);
when x"bb6" => lut_sig <= to_unsigned(integer(my_cos(2998)),16);
when x"bb7" => lut_sig <= to_unsigned(integer(my_cos(2999)),16);
when x"bb8" => lut_sig <= to_unsigned(integer(my_cos(3000)),16);
when x"bb9" => lut_sig <= to_unsigned(integer(my_cos(3001)),16);
when x"bba" => lut_sig <= to_unsigned(integer(my_cos(3002)),16);
when x"bbb" => lut_sig <= to_unsigned(integer(my_cos(3003)),16);
when x"bbc" => lut_sig <= to_unsigned(integer(my_cos(3004)),16);
when x"bbd" => lut_sig <= to_unsigned(integer(my_cos(3005)),16);
when x"bbe" => lut_sig <= to_unsigned(integer(my_cos(3006)),16);
when x"bbf" => lut_sig <= to_unsigned(integer(my_cos(3007)),16);
when x"bc0" => lut_sig <= to_unsigned(integer(my_cos(3008)),16);
when x"bc1" => lut_sig <= to_unsigned(integer(my_cos(3009)),16);
when x"bc2" => lut_sig <= to_unsigned(integer(my_cos(3010)),16);
when x"bc3" => lut_sig <= to_unsigned(integer(my_cos(3011)),16);
when x"bc4" => lut_sig <= to_unsigned(integer(my_cos(3012)),16);
when x"bc5" => lut_sig <= to_unsigned(integer(my_cos(3013)),16);
when x"bc6" => lut_sig <= to_unsigned(integer(my_cos(3014)),16);
when x"bc7" => lut_sig <= to_unsigned(integer(my_cos(3015)),16);
when x"bc8" => lut_sig <= to_unsigned(integer(my_cos(3016)),16);
when x"bc9" => lut_sig <= to_unsigned(integer(my_cos(3017)),16);
when x"bca" => lut_sig <= to_unsigned(integer(my_cos(3018)),16);
when x"bcb" => lut_sig <= to_unsigned(integer(my_cos(3019)),16);
when x"bcc" => lut_sig <= to_unsigned(integer(my_cos(3020)),16);
when x"bcd" => lut_sig <= to_unsigned(integer(my_cos(3021)),16);
when x"bce" => lut_sig <= to_unsigned(integer(my_cos(3022)),16);
when x"bcf" => lut_sig <= to_unsigned(integer(my_cos(3023)),16);
when x"bd0" => lut_sig <= to_unsigned(integer(my_cos(3024)),16);
when x"bd1" => lut_sig <= to_unsigned(integer(my_cos(3025)),16);
when x"bd2" => lut_sig <= to_unsigned(integer(my_cos(3026)),16);
when x"bd3" => lut_sig <= to_unsigned(integer(my_cos(3027)),16);
when x"bd4" => lut_sig <= to_unsigned(integer(my_cos(3028)),16);
when x"bd5" => lut_sig <= to_unsigned(integer(my_cos(3029)),16);
when x"bd6" => lut_sig <= to_unsigned(integer(my_cos(3030)),16);
when x"bd7" => lut_sig <= to_unsigned(integer(my_cos(3031)),16);
when x"bd8" => lut_sig <= to_unsigned(integer(my_cos(3032)),16);
when x"bd9" => lut_sig <= to_unsigned(integer(my_cos(3033)),16);
when x"bda" => lut_sig <= to_unsigned(integer(my_cos(3034)),16);
when x"bdb" => lut_sig <= to_unsigned(integer(my_cos(3035)),16);
when x"bdc" => lut_sig <= to_unsigned(integer(my_cos(3036)),16);
when x"bdd" => lut_sig <= to_unsigned(integer(my_cos(3037)),16);
when x"bde" => lut_sig <= to_unsigned(integer(my_cos(3038)),16);
when x"bdf" => lut_sig <= to_unsigned(integer(my_cos(3039)),16);
when x"be0" => lut_sig <= to_unsigned(integer(my_cos(3040)),16);
when x"be1" => lut_sig <= to_unsigned(integer(my_cos(3041)),16);
when x"be2" => lut_sig <= to_unsigned(integer(my_cos(3042)),16);
when x"be3" => lut_sig <= to_unsigned(integer(my_cos(3043)),16);
when x"be4" => lut_sig <= to_unsigned(integer(my_cos(3044)),16);
when x"be5" => lut_sig <= to_unsigned(integer(my_cos(3045)),16);
when x"be6" => lut_sig <= to_unsigned(integer(my_cos(3046)),16);
when x"be7" => lut_sig <= to_unsigned(integer(my_cos(3047)),16);
when x"be8" => lut_sig <= to_unsigned(integer(my_cos(3048)),16);
when x"be9" => lut_sig <= to_unsigned(integer(my_cos(3049)),16);
when x"bea" => lut_sig <= to_unsigned(integer(my_cos(3050)),16);
when x"beb" => lut_sig <= to_unsigned(integer(my_cos(3051)),16);
when x"bec" => lut_sig <= to_unsigned(integer(my_cos(3052)),16);
when x"bed" => lut_sig <= to_unsigned(integer(my_cos(3053)),16);
when x"bee" => lut_sig <= to_unsigned(integer(my_cos(3054)),16);
when x"bef" => lut_sig <= to_unsigned(integer(my_cos(3055)),16);
when x"bf0" => lut_sig <= to_unsigned(integer(my_cos(3056)),16);
when x"bf1" => lut_sig <= to_unsigned(integer(my_cos(3057)),16);
when x"bf2" => lut_sig <= to_unsigned(integer(my_cos(3058)),16);
when x"bf3" => lut_sig <= to_unsigned(integer(my_cos(3059)),16);
when x"bf4" => lut_sig <= to_unsigned(integer(my_cos(3060)),16);
when x"bf5" => lut_sig <= to_unsigned(integer(my_cos(3061)),16);
when x"bf6" => lut_sig <= to_unsigned(integer(my_cos(3062)),16);
when x"bf7" => lut_sig <= to_unsigned(integer(my_cos(3063)),16);
when x"bf8" => lut_sig <= to_unsigned(integer(my_cos(3064)),16);
when x"bf9" => lut_sig <= to_unsigned(integer(my_cos(3065)),16);
when x"bfa" => lut_sig <= to_unsigned(integer(my_cos(3066)),16);
when x"bfb" => lut_sig <= to_unsigned(integer(my_cos(3067)),16);
when x"bfc" => lut_sig <= to_unsigned(integer(my_cos(3068)),16);
when x"bfd" => lut_sig <= to_unsigned(integer(my_cos(3069)),16);
when x"bfe" => lut_sig <= to_unsigned(integer(my_cos(3070)),16);
when x"bff" => lut_sig <= to_unsigned(integer(my_cos(3071)),16);
when x"c00" => lut_sig <= to_unsigned(integer(my_cos(3072)),16);
when x"c01" => lut_sig <= to_unsigned(integer(my_cos(3073)),16);
when x"c02" => lut_sig <= to_unsigned(integer(my_cos(3074)),16);
when x"c03" => lut_sig <= to_unsigned(integer(my_cos(3075)),16);
when x"c04" => lut_sig <= to_unsigned(integer(my_cos(3076)),16);
when x"c05" => lut_sig <= to_unsigned(integer(my_cos(3077)),16);
when x"c06" => lut_sig <= to_unsigned(integer(my_cos(3078)),16);
when x"c07" => lut_sig <= to_unsigned(integer(my_cos(3079)),16);
when x"c08" => lut_sig <= to_unsigned(integer(my_cos(3080)),16);
when x"c09" => lut_sig <= to_unsigned(integer(my_cos(3081)),16);
when x"c0a" => lut_sig <= to_unsigned(integer(my_cos(3082)),16);
when x"c0b" => lut_sig <= to_unsigned(integer(my_cos(3083)),16);
when x"c0c" => lut_sig <= to_unsigned(integer(my_cos(3084)),16);
when x"c0d" => lut_sig <= to_unsigned(integer(my_cos(3085)),16);
when x"c0e" => lut_sig <= to_unsigned(integer(my_cos(3086)),16);
when x"c0f" => lut_sig <= to_unsigned(integer(my_cos(3087)),16);
when x"c10" => lut_sig <= to_unsigned(integer(my_cos(3088)),16);
when x"c11" => lut_sig <= to_unsigned(integer(my_cos(3089)),16);
when x"c12" => lut_sig <= to_unsigned(integer(my_cos(3090)),16);
when x"c13" => lut_sig <= to_unsigned(integer(my_cos(3091)),16);
when x"c14" => lut_sig <= to_unsigned(integer(my_cos(3092)),16);
when x"c15" => lut_sig <= to_unsigned(integer(my_cos(3093)),16);
when x"c16" => lut_sig <= to_unsigned(integer(my_cos(3094)),16);
when x"c17" => lut_sig <= to_unsigned(integer(my_cos(3095)),16);
when x"c18" => lut_sig <= to_unsigned(integer(my_cos(3096)),16);
when x"c19" => lut_sig <= to_unsigned(integer(my_cos(3097)),16);
when x"c1a" => lut_sig <= to_unsigned(integer(my_cos(3098)),16);
when x"c1b" => lut_sig <= to_unsigned(integer(my_cos(3099)),16);
when x"c1c" => lut_sig <= to_unsigned(integer(my_cos(3100)),16);
when x"c1d" => lut_sig <= to_unsigned(integer(my_cos(3101)),16);
when x"c1e" => lut_sig <= to_unsigned(integer(my_cos(3102)),16);
when x"c1f" => lut_sig <= to_unsigned(integer(my_cos(3103)),16);
when x"c20" => lut_sig <= to_unsigned(integer(my_cos(3104)),16);
when x"c21" => lut_sig <= to_unsigned(integer(my_cos(3105)),16);
when x"c22" => lut_sig <= to_unsigned(integer(my_cos(3106)),16);
when x"c23" => lut_sig <= to_unsigned(integer(my_cos(3107)),16);
when x"c24" => lut_sig <= to_unsigned(integer(my_cos(3108)),16);
when x"c25" => lut_sig <= to_unsigned(integer(my_cos(3109)),16);
when x"c26" => lut_sig <= to_unsigned(integer(my_cos(3110)),16);
when x"c27" => lut_sig <= to_unsigned(integer(my_cos(3111)),16);
when x"c28" => lut_sig <= to_unsigned(integer(my_cos(3112)),16);
when x"c29" => lut_sig <= to_unsigned(integer(my_cos(3113)),16);
when x"c2a" => lut_sig <= to_unsigned(integer(my_cos(3114)),16);
when x"c2b" => lut_sig <= to_unsigned(integer(my_cos(3115)),16);
when x"c2c" => lut_sig <= to_unsigned(integer(my_cos(3116)),16);
when x"c2d" => lut_sig <= to_unsigned(integer(my_cos(3117)),16);
when x"c2e" => lut_sig <= to_unsigned(integer(my_cos(3118)),16);
when x"c2f" => lut_sig <= to_unsigned(integer(my_cos(3119)),16);
when x"c30" => lut_sig <= to_unsigned(integer(my_cos(3120)),16);
when x"c31" => lut_sig <= to_unsigned(integer(my_cos(3121)),16);
when x"c32" => lut_sig <= to_unsigned(integer(my_cos(3122)),16);
when x"c33" => lut_sig <= to_unsigned(integer(my_cos(3123)),16);
when x"c34" => lut_sig <= to_unsigned(integer(my_cos(3124)),16);
when x"c35" => lut_sig <= to_unsigned(integer(my_cos(3125)),16);
when x"c36" => lut_sig <= to_unsigned(integer(my_cos(3126)),16);
when x"c37" => lut_sig <= to_unsigned(integer(my_cos(3127)),16);
when x"c38" => lut_sig <= to_unsigned(integer(my_cos(3128)),16);
when x"c39" => lut_sig <= to_unsigned(integer(my_cos(3129)),16);
when x"c3a" => lut_sig <= to_unsigned(integer(my_cos(3130)),16);
when x"c3b" => lut_sig <= to_unsigned(integer(my_cos(3131)),16);
when x"c3c" => lut_sig <= to_unsigned(integer(my_cos(3132)),16);
when x"c3d" => lut_sig <= to_unsigned(integer(my_cos(3133)),16);
when x"c3e" => lut_sig <= to_unsigned(integer(my_cos(3134)),16);
when x"c3f" => lut_sig <= to_unsigned(integer(my_cos(3135)),16);
when x"c40" => lut_sig <= to_unsigned(integer(my_cos(3136)),16);
when x"c41" => lut_sig <= to_unsigned(integer(my_cos(3137)),16);
when x"c42" => lut_sig <= to_unsigned(integer(my_cos(3138)),16);
when x"c43" => lut_sig <= to_unsigned(integer(my_cos(3139)),16);
when x"c44" => lut_sig <= to_unsigned(integer(my_cos(3140)),16);
when x"c45" => lut_sig <= to_unsigned(integer(my_cos(3141)),16);
when x"c46" => lut_sig <= to_unsigned(integer(my_cos(3142)),16);
when x"c47" => lut_sig <= to_unsigned(integer(my_cos(3143)),16);
when x"c48" => lut_sig <= to_unsigned(integer(my_cos(3144)),16);
when x"c49" => lut_sig <= to_unsigned(integer(my_cos(3145)),16);
when x"c4a" => lut_sig <= to_unsigned(integer(my_cos(3146)),16);
when x"c4b" => lut_sig <= to_unsigned(integer(my_cos(3147)),16);
when x"c4c" => lut_sig <= to_unsigned(integer(my_cos(3148)),16);
when x"c4d" => lut_sig <= to_unsigned(integer(my_cos(3149)),16);
when x"c4e" => lut_sig <= to_unsigned(integer(my_cos(3150)),16);
when x"c4f" => lut_sig <= to_unsigned(integer(my_cos(3151)),16);
when x"c50" => lut_sig <= to_unsigned(integer(my_cos(3152)),16);
when x"c51" => lut_sig <= to_unsigned(integer(my_cos(3153)),16);
when x"c52" => lut_sig <= to_unsigned(integer(my_cos(3154)),16);
when x"c53" => lut_sig <= to_unsigned(integer(my_cos(3155)),16);
when x"c54" => lut_sig <= to_unsigned(integer(my_cos(3156)),16);
when x"c55" => lut_sig <= to_unsigned(integer(my_cos(3157)),16);
when x"c56" => lut_sig <= to_unsigned(integer(my_cos(3158)),16);
when x"c57" => lut_sig <= to_unsigned(integer(my_cos(3159)),16);
when x"c58" => lut_sig <= to_unsigned(integer(my_cos(3160)),16);
when x"c59" => lut_sig <= to_unsigned(integer(my_cos(3161)),16);
when x"c5a" => lut_sig <= to_unsigned(integer(my_cos(3162)),16);
when x"c5b" => lut_sig <= to_unsigned(integer(my_cos(3163)),16);
when x"c5c" => lut_sig <= to_unsigned(integer(my_cos(3164)),16);
when x"c5d" => lut_sig <= to_unsigned(integer(my_cos(3165)),16);
when x"c5e" => lut_sig <= to_unsigned(integer(my_cos(3166)),16);
when x"c5f" => lut_sig <= to_unsigned(integer(my_cos(3167)),16);
when x"c60" => lut_sig <= to_unsigned(integer(my_cos(3168)),16);
when x"c61" => lut_sig <= to_unsigned(integer(my_cos(3169)),16);
when x"c62" => lut_sig <= to_unsigned(integer(my_cos(3170)),16);
when x"c63" => lut_sig <= to_unsigned(integer(my_cos(3171)),16);
when x"c64" => lut_sig <= to_unsigned(integer(my_cos(3172)),16);
when x"c65" => lut_sig <= to_unsigned(integer(my_cos(3173)),16);
when x"c66" => lut_sig <= to_unsigned(integer(my_cos(3174)),16);
when x"c67" => lut_sig <= to_unsigned(integer(my_cos(3175)),16);
when x"c68" => lut_sig <= to_unsigned(integer(my_cos(3176)),16);
when x"c69" => lut_sig <= to_unsigned(integer(my_cos(3177)),16);
when x"c6a" => lut_sig <= to_unsigned(integer(my_cos(3178)),16);
when x"c6b" => lut_sig <= to_unsigned(integer(my_cos(3179)),16);
when x"c6c" => lut_sig <= to_unsigned(integer(my_cos(3180)),16);
when x"c6d" => lut_sig <= to_unsigned(integer(my_cos(3181)),16);
when x"c6e" => lut_sig <= to_unsigned(integer(my_cos(3182)),16);
when x"c6f" => lut_sig <= to_unsigned(integer(my_cos(3183)),16);
when x"c70" => lut_sig <= to_unsigned(integer(my_cos(3184)),16);
when x"c71" => lut_sig <= to_unsigned(integer(my_cos(3185)),16);
when x"c72" => lut_sig <= to_unsigned(integer(my_cos(3186)),16);
when x"c73" => lut_sig <= to_unsigned(integer(my_cos(3187)),16);
when x"c74" => lut_sig <= to_unsigned(integer(my_cos(3188)),16);
when x"c75" => lut_sig <= to_unsigned(integer(my_cos(3189)),16);
when x"c76" => lut_sig <= to_unsigned(integer(my_cos(3190)),16);
when x"c77" => lut_sig <= to_unsigned(integer(my_cos(3191)),16);
when x"c78" => lut_sig <= to_unsigned(integer(my_cos(3192)),16);
when x"c79" => lut_sig <= to_unsigned(integer(my_cos(3193)),16);
when x"c7a" => lut_sig <= to_unsigned(integer(my_cos(3194)),16);
when x"c7b" => lut_sig <= to_unsigned(integer(my_cos(3195)),16);
when x"c7c" => lut_sig <= to_unsigned(integer(my_cos(3196)),16);
when x"c7d" => lut_sig <= to_unsigned(integer(my_cos(3197)),16);
when x"c7e" => lut_sig <= to_unsigned(integer(my_cos(3198)),16);
when x"c7f" => lut_sig <= to_unsigned(integer(my_cos(3199)),16);
when x"c80" => lut_sig <= to_unsigned(integer(my_cos(3200)),16);
when x"c81" => lut_sig <= to_unsigned(integer(my_cos(3201)),16);
when x"c82" => lut_sig <= to_unsigned(integer(my_cos(3202)),16);
when x"c83" => lut_sig <= to_unsigned(integer(my_cos(3203)),16);
when x"c84" => lut_sig <= to_unsigned(integer(my_cos(3204)),16);
when x"c85" => lut_sig <= to_unsigned(integer(my_cos(3205)),16);
when x"c86" => lut_sig <= to_unsigned(integer(my_cos(3206)),16);
when x"c87" => lut_sig <= to_unsigned(integer(my_cos(3207)),16);
when x"c88" => lut_sig <= to_unsigned(integer(my_cos(3208)),16);
when x"c89" => lut_sig <= to_unsigned(integer(my_cos(3209)),16);
when x"c8a" => lut_sig <= to_unsigned(integer(my_cos(3210)),16);
when x"c8b" => lut_sig <= to_unsigned(integer(my_cos(3211)),16);
when x"c8c" => lut_sig <= to_unsigned(integer(my_cos(3212)),16);
when x"c8d" => lut_sig <= to_unsigned(integer(my_cos(3213)),16);
when x"c8e" => lut_sig <= to_unsigned(integer(my_cos(3214)),16);
when x"c8f" => lut_sig <= to_unsigned(integer(my_cos(3215)),16);
when x"c90" => lut_sig <= to_unsigned(integer(my_cos(3216)),16);
when x"c91" => lut_sig <= to_unsigned(integer(my_cos(3217)),16);
when x"c92" => lut_sig <= to_unsigned(integer(my_cos(3218)),16);
when x"c93" => lut_sig <= to_unsigned(integer(my_cos(3219)),16);
when x"c94" => lut_sig <= to_unsigned(integer(my_cos(3220)),16);
when x"c95" => lut_sig <= to_unsigned(integer(my_cos(3221)),16);
when x"c96" => lut_sig <= to_unsigned(integer(my_cos(3222)),16);
when x"c97" => lut_sig <= to_unsigned(integer(my_cos(3223)),16);
when x"c98" => lut_sig <= to_unsigned(integer(my_cos(3224)),16);
when x"c99" => lut_sig <= to_unsigned(integer(my_cos(3225)),16);
when x"c9a" => lut_sig <= to_unsigned(integer(my_cos(3226)),16);
when x"c9b" => lut_sig <= to_unsigned(integer(my_cos(3227)),16);
when x"c9c" => lut_sig <= to_unsigned(integer(my_cos(3228)),16);
when x"c9d" => lut_sig <= to_unsigned(integer(my_cos(3229)),16);
when x"c9e" => lut_sig <= to_unsigned(integer(my_cos(3230)),16);
when x"c9f" => lut_sig <= to_unsigned(integer(my_cos(3231)),16);
when x"ca0" => lut_sig <= to_unsigned(integer(my_cos(3232)),16);
when x"ca1" => lut_sig <= to_unsigned(integer(my_cos(3233)),16);
when x"ca2" => lut_sig <= to_unsigned(integer(my_cos(3234)),16);
when x"ca3" => lut_sig <= to_unsigned(integer(my_cos(3235)),16);
when x"ca4" => lut_sig <= to_unsigned(integer(my_cos(3236)),16);
when x"ca5" => lut_sig <= to_unsigned(integer(my_cos(3237)),16);
when x"ca6" => lut_sig <= to_unsigned(integer(my_cos(3238)),16);
when x"ca7" => lut_sig <= to_unsigned(integer(my_cos(3239)),16);
when x"ca8" => lut_sig <= to_unsigned(integer(my_cos(3240)),16);
when x"ca9" => lut_sig <= to_unsigned(integer(my_cos(3241)),16);
when x"caa" => lut_sig <= to_unsigned(integer(my_cos(3242)),16);
when x"cab" => lut_sig <= to_unsigned(integer(my_cos(3243)),16);
when x"cac" => lut_sig <= to_unsigned(integer(my_cos(3244)),16);
when x"cad" => lut_sig <= to_unsigned(integer(my_cos(3245)),16);
when x"cae" => lut_sig <= to_unsigned(integer(my_cos(3246)),16);
when x"caf" => lut_sig <= to_unsigned(integer(my_cos(3247)),16);
when x"cb0" => lut_sig <= to_unsigned(integer(my_cos(3248)),16);
when x"cb1" => lut_sig <= to_unsigned(integer(my_cos(3249)),16);
when x"cb2" => lut_sig <= to_unsigned(integer(my_cos(3250)),16);
when x"cb3" => lut_sig <= to_unsigned(integer(my_cos(3251)),16);
when x"cb4" => lut_sig <= to_unsigned(integer(my_cos(3252)),16);
when x"cb5" => lut_sig <= to_unsigned(integer(my_cos(3253)),16);
when x"cb6" => lut_sig <= to_unsigned(integer(my_cos(3254)),16);
when x"cb7" => lut_sig <= to_unsigned(integer(my_cos(3255)),16);
when x"cb8" => lut_sig <= to_unsigned(integer(my_cos(3256)),16);
when x"cb9" => lut_sig <= to_unsigned(integer(my_cos(3257)),16);
when x"cba" => lut_sig <= to_unsigned(integer(my_cos(3258)),16);
when x"cbb" => lut_sig <= to_unsigned(integer(my_cos(3259)),16);
when x"cbc" => lut_sig <= to_unsigned(integer(my_cos(3260)),16);
when x"cbd" => lut_sig <= to_unsigned(integer(my_cos(3261)),16);
when x"cbe" => lut_sig <= to_unsigned(integer(my_cos(3262)),16);
when x"cbf" => lut_sig <= to_unsigned(integer(my_cos(3263)),16);
when x"cc0" => lut_sig <= to_unsigned(integer(my_cos(3264)),16);
when x"cc1" => lut_sig <= to_unsigned(integer(my_cos(3265)),16);
when x"cc2" => lut_sig <= to_unsigned(integer(my_cos(3266)),16);
when x"cc3" => lut_sig <= to_unsigned(integer(my_cos(3267)),16);
when x"cc4" => lut_sig <= to_unsigned(integer(my_cos(3268)),16);
when x"cc5" => lut_sig <= to_unsigned(integer(my_cos(3269)),16);
when x"cc6" => lut_sig <= to_unsigned(integer(my_cos(3270)),16);
when x"cc7" => lut_sig <= to_unsigned(integer(my_cos(3271)),16);
when x"cc8" => lut_sig <= to_unsigned(integer(my_cos(3272)),16);
when x"cc9" => lut_sig <= to_unsigned(integer(my_cos(3273)),16);
when x"cca" => lut_sig <= to_unsigned(integer(my_cos(3274)),16);
when x"ccb" => lut_sig <= to_unsigned(integer(my_cos(3275)),16);
when x"ccc" => lut_sig <= to_unsigned(integer(my_cos(3276)),16);
when x"ccd" => lut_sig <= to_unsigned(integer(my_cos(3277)),16);
when x"cce" => lut_sig <= to_unsigned(integer(my_cos(3278)),16);
when x"ccf" => lut_sig <= to_unsigned(integer(my_cos(3279)),16);
when x"cd0" => lut_sig <= to_unsigned(integer(my_cos(3280)),16);
when x"cd1" => lut_sig <= to_unsigned(integer(my_cos(3281)),16);
when x"cd2" => lut_sig <= to_unsigned(integer(my_cos(3282)),16);
when x"cd3" => lut_sig <= to_unsigned(integer(my_cos(3283)),16);
when x"cd4" => lut_sig <= to_unsigned(integer(my_cos(3284)),16);
when x"cd5" => lut_sig <= to_unsigned(integer(my_cos(3285)),16);
when x"cd6" => lut_sig <= to_unsigned(integer(my_cos(3286)),16);
when x"cd7" => lut_sig <= to_unsigned(integer(my_cos(3287)),16);
when x"cd8" => lut_sig <= to_unsigned(integer(my_cos(3288)),16);
when x"cd9" => lut_sig <= to_unsigned(integer(my_cos(3289)),16);
when x"cda" => lut_sig <= to_unsigned(integer(my_cos(3290)),16);
when x"cdb" => lut_sig <= to_unsigned(integer(my_cos(3291)),16);
when x"cdc" => lut_sig <= to_unsigned(integer(my_cos(3292)),16);
when x"cdd" => lut_sig <= to_unsigned(integer(my_cos(3293)),16);
when x"cde" => lut_sig <= to_unsigned(integer(my_cos(3294)),16);
when x"cdf" => lut_sig <= to_unsigned(integer(my_cos(3295)),16);
when x"ce0" => lut_sig <= to_unsigned(integer(my_cos(3296)),16);
when x"ce1" => lut_sig <= to_unsigned(integer(my_cos(3297)),16);
when x"ce2" => lut_sig <= to_unsigned(integer(my_cos(3298)),16);
when x"ce3" => lut_sig <= to_unsigned(integer(my_cos(3299)),16);
when x"ce4" => lut_sig <= to_unsigned(integer(my_cos(3300)),16);
when x"ce5" => lut_sig <= to_unsigned(integer(my_cos(3301)),16);
when x"ce6" => lut_sig <= to_unsigned(integer(my_cos(3302)),16);
when x"ce7" => lut_sig <= to_unsigned(integer(my_cos(3303)),16);
when x"ce8" => lut_sig <= to_unsigned(integer(my_cos(3304)),16);
when x"ce9" => lut_sig <= to_unsigned(integer(my_cos(3305)),16);
when x"cea" => lut_sig <= to_unsigned(integer(my_cos(3306)),16);
when x"ceb" => lut_sig <= to_unsigned(integer(my_cos(3307)),16);
when x"cec" => lut_sig <= to_unsigned(integer(my_cos(3308)),16);
when x"ced" => lut_sig <= to_unsigned(integer(my_cos(3309)),16);
when x"cee" => lut_sig <= to_unsigned(integer(my_cos(3310)),16);
when x"cef" => lut_sig <= to_unsigned(integer(my_cos(3311)),16);
when x"cf0" => lut_sig <= to_unsigned(integer(my_cos(3312)),16);
when x"cf1" => lut_sig <= to_unsigned(integer(my_cos(3313)),16);
when x"cf2" => lut_sig <= to_unsigned(integer(my_cos(3314)),16);
when x"cf3" => lut_sig <= to_unsigned(integer(my_cos(3315)),16);
when x"cf4" => lut_sig <= to_unsigned(integer(my_cos(3316)),16);
when x"cf5" => lut_sig <= to_unsigned(integer(my_cos(3317)),16);
when x"cf6" => lut_sig <= to_unsigned(integer(my_cos(3318)),16);
when x"cf7" => lut_sig <= to_unsigned(integer(my_cos(3319)),16);
when x"cf8" => lut_sig <= to_unsigned(integer(my_cos(3320)),16);
when x"cf9" => lut_sig <= to_unsigned(integer(my_cos(3321)),16);
when x"cfa" => lut_sig <= to_unsigned(integer(my_cos(3322)),16);
when x"cfb" => lut_sig <= to_unsigned(integer(my_cos(3323)),16);
when x"cfc" => lut_sig <= to_unsigned(integer(my_cos(3324)),16);
when x"cfd" => lut_sig <= to_unsigned(integer(my_cos(3325)),16);
when x"cfe" => lut_sig <= to_unsigned(integer(my_cos(3326)),16);
when x"cff" => lut_sig <= to_unsigned(integer(my_cos(3327)),16);
when x"d00" => lut_sig <= to_unsigned(integer(my_cos(3328)),16);
when x"d01" => lut_sig <= to_unsigned(integer(my_cos(3329)),16);
when x"d02" => lut_sig <= to_unsigned(integer(my_cos(3330)),16);
when x"d03" => lut_sig <= to_unsigned(integer(my_cos(3331)),16);
when x"d04" => lut_sig <= to_unsigned(integer(my_cos(3332)),16);
when x"d05" => lut_sig <= to_unsigned(integer(my_cos(3333)),16);
when x"d06" => lut_sig <= to_unsigned(integer(my_cos(3334)),16);
when x"d07" => lut_sig <= to_unsigned(integer(my_cos(3335)),16);
when x"d08" => lut_sig <= to_unsigned(integer(my_cos(3336)),16);
when x"d09" => lut_sig <= to_unsigned(integer(my_cos(3337)),16);
when x"d0a" => lut_sig <= to_unsigned(integer(my_cos(3338)),16);
when x"d0b" => lut_sig <= to_unsigned(integer(my_cos(3339)),16);
when x"d0c" => lut_sig <= to_unsigned(integer(my_cos(3340)),16);
when x"d0d" => lut_sig <= to_unsigned(integer(my_cos(3341)),16);
when x"d0e" => lut_sig <= to_unsigned(integer(my_cos(3342)),16);
when x"d0f" => lut_sig <= to_unsigned(integer(my_cos(3343)),16);
when x"d10" => lut_sig <= to_unsigned(integer(my_cos(3344)),16);
when x"d11" => lut_sig <= to_unsigned(integer(my_cos(3345)),16);
when x"d12" => lut_sig <= to_unsigned(integer(my_cos(3346)),16);
when x"d13" => lut_sig <= to_unsigned(integer(my_cos(3347)),16);
when x"d14" => lut_sig <= to_unsigned(integer(my_cos(3348)),16);
when x"d15" => lut_sig <= to_unsigned(integer(my_cos(3349)),16);
when x"d16" => lut_sig <= to_unsigned(integer(my_cos(3350)),16);
when x"d17" => lut_sig <= to_unsigned(integer(my_cos(3351)),16);
when x"d18" => lut_sig <= to_unsigned(integer(my_cos(3352)),16);
when x"d19" => lut_sig <= to_unsigned(integer(my_cos(3353)),16);
when x"d1a" => lut_sig <= to_unsigned(integer(my_cos(3354)),16);
when x"d1b" => lut_sig <= to_unsigned(integer(my_cos(3355)),16);
when x"d1c" => lut_sig <= to_unsigned(integer(my_cos(3356)),16);
when x"d1d" => lut_sig <= to_unsigned(integer(my_cos(3357)),16);
when x"d1e" => lut_sig <= to_unsigned(integer(my_cos(3358)),16);
when x"d1f" => lut_sig <= to_unsigned(integer(my_cos(3359)),16);
when x"d20" => lut_sig <= to_unsigned(integer(my_cos(3360)),16);
when x"d21" => lut_sig <= to_unsigned(integer(my_cos(3361)),16);
when x"d22" => lut_sig <= to_unsigned(integer(my_cos(3362)),16);
when x"d23" => lut_sig <= to_unsigned(integer(my_cos(3363)),16);
when x"d24" => lut_sig <= to_unsigned(integer(my_cos(3364)),16);
when x"d25" => lut_sig <= to_unsigned(integer(my_cos(3365)),16);
when x"d26" => lut_sig <= to_unsigned(integer(my_cos(3366)),16);
when x"d27" => lut_sig <= to_unsigned(integer(my_cos(3367)),16);
when x"d28" => lut_sig <= to_unsigned(integer(my_cos(3368)),16);
when x"d29" => lut_sig <= to_unsigned(integer(my_cos(3369)),16);
when x"d2a" => lut_sig <= to_unsigned(integer(my_cos(3370)),16);
when x"d2b" => lut_sig <= to_unsigned(integer(my_cos(3371)),16);
when x"d2c" => lut_sig <= to_unsigned(integer(my_cos(3372)),16);
when x"d2d" => lut_sig <= to_unsigned(integer(my_cos(3373)),16);
when x"d2e" => lut_sig <= to_unsigned(integer(my_cos(3374)),16);
when x"d2f" => lut_sig <= to_unsigned(integer(my_cos(3375)),16);
when x"d30" => lut_sig <= to_unsigned(integer(my_cos(3376)),16);
when x"d31" => lut_sig <= to_unsigned(integer(my_cos(3377)),16);
when x"d32" => lut_sig <= to_unsigned(integer(my_cos(3378)),16);
when x"d33" => lut_sig <= to_unsigned(integer(my_cos(3379)),16);
when x"d34" => lut_sig <= to_unsigned(integer(my_cos(3380)),16);
when x"d35" => lut_sig <= to_unsigned(integer(my_cos(3381)),16);
when x"d36" => lut_sig <= to_unsigned(integer(my_cos(3382)),16);
when x"d37" => lut_sig <= to_unsigned(integer(my_cos(3383)),16);
when x"d38" => lut_sig <= to_unsigned(integer(my_cos(3384)),16);
when x"d39" => lut_sig <= to_unsigned(integer(my_cos(3385)),16);
when x"d3a" => lut_sig <= to_unsigned(integer(my_cos(3386)),16);
when x"d3b" => lut_sig <= to_unsigned(integer(my_cos(3387)),16);
when x"d3c" => lut_sig <= to_unsigned(integer(my_cos(3388)),16);
when x"d3d" => lut_sig <= to_unsigned(integer(my_cos(3389)),16);
when x"d3e" => lut_sig <= to_unsigned(integer(my_cos(3390)),16);
when x"d3f" => lut_sig <= to_unsigned(integer(my_cos(3391)),16);
when x"d40" => lut_sig <= to_unsigned(integer(my_cos(3392)),16);
when x"d41" => lut_sig <= to_unsigned(integer(my_cos(3393)),16);
when x"d42" => lut_sig <= to_unsigned(integer(my_cos(3394)),16);
when x"d43" => lut_sig <= to_unsigned(integer(my_cos(3395)),16);
when x"d44" => lut_sig <= to_unsigned(integer(my_cos(3396)),16);
when x"d45" => lut_sig <= to_unsigned(integer(my_cos(3397)),16);
when x"d46" => lut_sig <= to_unsigned(integer(my_cos(3398)),16);
when x"d47" => lut_sig <= to_unsigned(integer(my_cos(3399)),16);
when x"d48" => lut_sig <= to_unsigned(integer(my_cos(3400)),16);
when x"d49" => lut_sig <= to_unsigned(integer(my_cos(3401)),16);
when x"d4a" => lut_sig <= to_unsigned(integer(my_cos(3402)),16);
when x"d4b" => lut_sig <= to_unsigned(integer(my_cos(3403)),16);
when x"d4c" => lut_sig <= to_unsigned(integer(my_cos(3404)),16);
when x"d4d" => lut_sig <= to_unsigned(integer(my_cos(3405)),16);
when x"d4e" => lut_sig <= to_unsigned(integer(my_cos(3406)),16);
when x"d4f" => lut_sig <= to_unsigned(integer(my_cos(3407)),16);
when x"d50" => lut_sig <= to_unsigned(integer(my_cos(3408)),16);
when x"d51" => lut_sig <= to_unsigned(integer(my_cos(3409)),16);
when x"d52" => lut_sig <= to_unsigned(integer(my_cos(3410)),16);
when x"d53" => lut_sig <= to_unsigned(integer(my_cos(3411)),16);
when x"d54" => lut_sig <= to_unsigned(integer(my_cos(3412)),16);
when x"d55" => lut_sig <= to_unsigned(integer(my_cos(3413)),16);
when x"d56" => lut_sig <= to_unsigned(integer(my_cos(3414)),16);
when x"d57" => lut_sig <= to_unsigned(integer(my_cos(3415)),16);
when x"d58" => lut_sig <= to_unsigned(integer(my_cos(3416)),16);
when x"d59" => lut_sig <= to_unsigned(integer(my_cos(3417)),16);
when x"d5a" => lut_sig <= to_unsigned(integer(my_cos(3418)),16);
when x"d5b" => lut_sig <= to_unsigned(integer(my_cos(3419)),16);
when x"d5c" => lut_sig <= to_unsigned(integer(my_cos(3420)),16);
when x"d5d" => lut_sig <= to_unsigned(integer(my_cos(3421)),16);
when x"d5e" => lut_sig <= to_unsigned(integer(my_cos(3422)),16);
when x"d5f" => lut_sig <= to_unsigned(integer(my_cos(3423)),16);
when x"d60" => lut_sig <= to_unsigned(integer(my_cos(3424)),16);
when x"d61" => lut_sig <= to_unsigned(integer(my_cos(3425)),16);
when x"d62" => lut_sig <= to_unsigned(integer(my_cos(3426)),16);
when x"d63" => lut_sig <= to_unsigned(integer(my_cos(3427)),16);
when x"d64" => lut_sig <= to_unsigned(integer(my_cos(3428)),16);
when x"d65" => lut_sig <= to_unsigned(integer(my_cos(3429)),16);
when x"d66" => lut_sig <= to_unsigned(integer(my_cos(3430)),16);
when x"d67" => lut_sig <= to_unsigned(integer(my_cos(3431)),16);
when x"d68" => lut_sig <= to_unsigned(integer(my_cos(3432)),16);
when x"d69" => lut_sig <= to_unsigned(integer(my_cos(3433)),16);
when x"d6a" => lut_sig <= to_unsigned(integer(my_cos(3434)),16);
when x"d6b" => lut_sig <= to_unsigned(integer(my_cos(3435)),16);
when x"d6c" => lut_sig <= to_unsigned(integer(my_cos(3436)),16);
when x"d6d" => lut_sig <= to_unsigned(integer(my_cos(3437)),16);
when x"d6e" => lut_sig <= to_unsigned(integer(my_cos(3438)),16);
when x"d6f" => lut_sig <= to_unsigned(integer(my_cos(3439)),16);
when x"d70" => lut_sig <= to_unsigned(integer(my_cos(3440)),16);
when x"d71" => lut_sig <= to_unsigned(integer(my_cos(3441)),16);
when x"d72" => lut_sig <= to_unsigned(integer(my_cos(3442)),16);
when x"d73" => lut_sig <= to_unsigned(integer(my_cos(3443)),16);
when x"d74" => lut_sig <= to_unsigned(integer(my_cos(3444)),16);
when x"d75" => lut_sig <= to_unsigned(integer(my_cos(3445)),16);
when x"d76" => lut_sig <= to_unsigned(integer(my_cos(3446)),16);
when x"d77" => lut_sig <= to_unsigned(integer(my_cos(3447)),16);
when x"d78" => lut_sig <= to_unsigned(integer(my_cos(3448)),16);
when x"d79" => lut_sig <= to_unsigned(integer(my_cos(3449)),16);
when x"d7a" => lut_sig <= to_unsigned(integer(my_cos(3450)),16);
when x"d7b" => lut_sig <= to_unsigned(integer(my_cos(3451)),16);
when x"d7c" => lut_sig <= to_unsigned(integer(my_cos(3452)),16);
when x"d7d" => lut_sig <= to_unsigned(integer(my_cos(3453)),16);
when x"d7e" => lut_sig <= to_unsigned(integer(my_cos(3454)),16);
when x"d7f" => lut_sig <= to_unsigned(integer(my_cos(3455)),16);
when x"d80" => lut_sig <= to_unsigned(integer(my_cos(3456)),16);
when x"d81" => lut_sig <= to_unsigned(integer(my_cos(3457)),16);
when x"d82" => lut_sig <= to_unsigned(integer(my_cos(3458)),16);
when x"d83" => lut_sig <= to_unsigned(integer(my_cos(3459)),16);
when x"d84" => lut_sig <= to_unsigned(integer(my_cos(3460)),16);
when x"d85" => lut_sig <= to_unsigned(integer(my_cos(3461)),16);
when x"d86" => lut_sig <= to_unsigned(integer(my_cos(3462)),16);
when x"d87" => lut_sig <= to_unsigned(integer(my_cos(3463)),16);
when x"d88" => lut_sig <= to_unsigned(integer(my_cos(3464)),16);
when x"d89" => lut_sig <= to_unsigned(integer(my_cos(3465)),16);
when x"d8a" => lut_sig <= to_unsigned(integer(my_cos(3466)),16);
when x"d8b" => lut_sig <= to_unsigned(integer(my_cos(3467)),16);
when x"d8c" => lut_sig <= to_unsigned(integer(my_cos(3468)),16);
when x"d8d" => lut_sig <= to_unsigned(integer(my_cos(3469)),16);
when x"d8e" => lut_sig <= to_unsigned(integer(my_cos(3470)),16);
when x"d8f" => lut_sig <= to_unsigned(integer(my_cos(3471)),16);
when x"d90" => lut_sig <= to_unsigned(integer(my_cos(3472)),16);
when x"d91" => lut_sig <= to_unsigned(integer(my_cos(3473)),16);
when x"d92" => lut_sig <= to_unsigned(integer(my_cos(3474)),16);
when x"d93" => lut_sig <= to_unsigned(integer(my_cos(3475)),16);
when x"d94" => lut_sig <= to_unsigned(integer(my_cos(3476)),16);
when x"d95" => lut_sig <= to_unsigned(integer(my_cos(3477)),16);
when x"d96" => lut_sig <= to_unsigned(integer(my_cos(3478)),16);
when x"d97" => lut_sig <= to_unsigned(integer(my_cos(3479)),16);
when x"d98" => lut_sig <= to_unsigned(integer(my_cos(3480)),16);
when x"d99" => lut_sig <= to_unsigned(integer(my_cos(3481)),16);
when x"d9a" => lut_sig <= to_unsigned(integer(my_cos(3482)),16);
when x"d9b" => lut_sig <= to_unsigned(integer(my_cos(3483)),16);
when x"d9c" => lut_sig <= to_unsigned(integer(my_cos(3484)),16);
when x"d9d" => lut_sig <= to_unsigned(integer(my_cos(3485)),16);
when x"d9e" => lut_sig <= to_unsigned(integer(my_cos(3486)),16);
when x"d9f" => lut_sig <= to_unsigned(integer(my_cos(3487)),16);
when x"da0" => lut_sig <= to_unsigned(integer(my_cos(3488)),16);
when x"da1" => lut_sig <= to_unsigned(integer(my_cos(3489)),16);
when x"da2" => lut_sig <= to_unsigned(integer(my_cos(3490)),16);
when x"da3" => lut_sig <= to_unsigned(integer(my_cos(3491)),16);
when x"da4" => lut_sig <= to_unsigned(integer(my_cos(3492)),16);
when x"da5" => lut_sig <= to_unsigned(integer(my_cos(3493)),16);
when x"da6" => lut_sig <= to_unsigned(integer(my_cos(3494)),16);
when x"da7" => lut_sig <= to_unsigned(integer(my_cos(3495)),16);
when x"da8" => lut_sig <= to_unsigned(integer(my_cos(3496)),16);
when x"da9" => lut_sig <= to_unsigned(integer(my_cos(3497)),16);
when x"daa" => lut_sig <= to_unsigned(integer(my_cos(3498)),16);
when x"dab" => lut_sig <= to_unsigned(integer(my_cos(3499)),16);
when x"dac" => lut_sig <= to_unsigned(integer(my_cos(3500)),16);
when x"dad" => lut_sig <= to_unsigned(integer(my_cos(3501)),16);
when x"dae" => lut_sig <= to_unsigned(integer(my_cos(3502)),16);
when x"daf" => lut_sig <= to_unsigned(integer(my_cos(3503)),16);
when x"db0" => lut_sig <= to_unsigned(integer(my_cos(3504)),16);
when x"db1" => lut_sig <= to_unsigned(integer(my_cos(3505)),16);
when x"db2" => lut_sig <= to_unsigned(integer(my_cos(3506)),16);
when x"db3" => lut_sig <= to_unsigned(integer(my_cos(3507)),16);
when x"db4" => lut_sig <= to_unsigned(integer(my_cos(3508)),16);
when x"db5" => lut_sig <= to_unsigned(integer(my_cos(3509)),16);
when x"db6" => lut_sig <= to_unsigned(integer(my_cos(3510)),16);
when x"db7" => lut_sig <= to_unsigned(integer(my_cos(3511)),16);
when x"db8" => lut_sig <= to_unsigned(integer(my_cos(3512)),16);
when x"db9" => lut_sig <= to_unsigned(integer(my_cos(3513)),16);
when x"dba" => lut_sig <= to_unsigned(integer(my_cos(3514)),16);
when x"dbb" => lut_sig <= to_unsigned(integer(my_cos(3515)),16);
when x"dbc" => lut_sig <= to_unsigned(integer(my_cos(3516)),16);
when x"dbd" => lut_sig <= to_unsigned(integer(my_cos(3517)),16);
when x"dbe" => lut_sig <= to_unsigned(integer(my_cos(3518)),16);
when x"dbf" => lut_sig <= to_unsigned(integer(my_cos(3519)),16);
when x"dc0" => lut_sig <= to_unsigned(integer(my_cos(3520)),16);
when x"dc1" => lut_sig <= to_unsigned(integer(my_cos(3521)),16);
when x"dc2" => lut_sig <= to_unsigned(integer(my_cos(3522)),16);
when x"dc3" => lut_sig <= to_unsigned(integer(my_cos(3523)),16);
when x"dc4" => lut_sig <= to_unsigned(integer(my_cos(3524)),16);
when x"dc5" => lut_sig <= to_unsigned(integer(my_cos(3525)),16);
when x"dc6" => lut_sig <= to_unsigned(integer(my_cos(3526)),16);
when x"dc7" => lut_sig <= to_unsigned(integer(my_cos(3527)),16);
when x"dc8" => lut_sig <= to_unsigned(integer(my_cos(3528)),16);
when x"dc9" => lut_sig <= to_unsigned(integer(my_cos(3529)),16);
when x"dca" => lut_sig <= to_unsigned(integer(my_cos(3530)),16);
when x"dcb" => lut_sig <= to_unsigned(integer(my_cos(3531)),16);
when x"dcc" => lut_sig <= to_unsigned(integer(my_cos(3532)),16);
when x"dcd" => lut_sig <= to_unsigned(integer(my_cos(3533)),16);
when x"dce" => lut_sig <= to_unsigned(integer(my_cos(3534)),16);
when x"dcf" => lut_sig <= to_unsigned(integer(my_cos(3535)),16);
when x"dd0" => lut_sig <= to_unsigned(integer(my_cos(3536)),16);
when x"dd1" => lut_sig <= to_unsigned(integer(my_cos(3537)),16);
when x"dd2" => lut_sig <= to_unsigned(integer(my_cos(3538)),16);
when x"dd3" => lut_sig <= to_unsigned(integer(my_cos(3539)),16);
when x"dd4" => lut_sig <= to_unsigned(integer(my_cos(3540)),16);
when x"dd5" => lut_sig <= to_unsigned(integer(my_cos(3541)),16);
when x"dd6" => lut_sig <= to_unsigned(integer(my_cos(3542)),16);
when x"dd7" => lut_sig <= to_unsigned(integer(my_cos(3543)),16);
when x"dd8" => lut_sig <= to_unsigned(integer(my_cos(3544)),16);
when x"dd9" => lut_sig <= to_unsigned(integer(my_cos(3545)),16);
when x"dda" => lut_sig <= to_unsigned(integer(my_cos(3546)),16);
when x"ddb" => lut_sig <= to_unsigned(integer(my_cos(3547)),16);
when x"ddc" => lut_sig <= to_unsigned(integer(my_cos(3548)),16);
when x"ddd" => lut_sig <= to_unsigned(integer(my_cos(3549)),16);
when x"dde" => lut_sig <= to_unsigned(integer(my_cos(3550)),16);
when x"ddf" => lut_sig <= to_unsigned(integer(my_cos(3551)),16);
when x"de0" => lut_sig <= to_unsigned(integer(my_cos(3552)),16);
when x"de1" => lut_sig <= to_unsigned(integer(my_cos(3553)),16);
when x"de2" => lut_sig <= to_unsigned(integer(my_cos(3554)),16);
when x"de3" => lut_sig <= to_unsigned(integer(my_cos(3555)),16);
when x"de4" => lut_sig <= to_unsigned(integer(my_cos(3556)),16);
when x"de5" => lut_sig <= to_unsigned(integer(my_cos(3557)),16);
when x"de6" => lut_sig <= to_unsigned(integer(my_cos(3558)),16);
when x"de7" => lut_sig <= to_unsigned(integer(my_cos(3559)),16);
when x"de8" => lut_sig <= to_unsigned(integer(my_cos(3560)),16);
when x"de9" => lut_sig <= to_unsigned(integer(my_cos(3561)),16);
when x"dea" => lut_sig <= to_unsigned(integer(my_cos(3562)),16);
when x"deb" => lut_sig <= to_unsigned(integer(my_cos(3563)),16);
when x"dec" => lut_sig <= to_unsigned(integer(my_cos(3564)),16);
when x"ded" => lut_sig <= to_unsigned(integer(my_cos(3565)),16);
when x"dee" => lut_sig <= to_unsigned(integer(my_cos(3566)),16);
when x"def" => lut_sig <= to_unsigned(integer(my_cos(3567)),16);
when x"df0" => lut_sig <= to_unsigned(integer(my_cos(3568)),16);
when x"df1" => lut_sig <= to_unsigned(integer(my_cos(3569)),16);
when x"df2" => lut_sig <= to_unsigned(integer(my_cos(3570)),16);
when x"df3" => lut_sig <= to_unsigned(integer(my_cos(3571)),16);
when x"df4" => lut_sig <= to_unsigned(integer(my_cos(3572)),16);
when x"df5" => lut_sig <= to_unsigned(integer(my_cos(3573)),16);
when x"df6" => lut_sig <= to_unsigned(integer(my_cos(3574)),16);
when x"df7" => lut_sig <= to_unsigned(integer(my_cos(3575)),16);
when x"df8" => lut_sig <= to_unsigned(integer(my_cos(3576)),16);
when x"df9" => lut_sig <= to_unsigned(integer(my_cos(3577)),16);
when x"dfa" => lut_sig <= to_unsigned(integer(my_cos(3578)),16);
when x"dfb" => lut_sig <= to_unsigned(integer(my_cos(3579)),16);
when x"dfc" => lut_sig <= to_unsigned(integer(my_cos(3580)),16);
when x"dfd" => lut_sig <= to_unsigned(integer(my_cos(3581)),16);
when x"dfe" => lut_sig <= to_unsigned(integer(my_cos(3582)),16);
when x"dff" => lut_sig <= to_unsigned(integer(my_cos(3583)),16);
when x"e00" => lut_sig <= to_unsigned(integer(my_cos(3584)),16);
when x"e01" => lut_sig <= to_unsigned(integer(my_cos(3585)),16);
when x"e02" => lut_sig <= to_unsigned(integer(my_cos(3586)),16);
when x"e03" => lut_sig <= to_unsigned(integer(my_cos(3587)),16);
when x"e04" => lut_sig <= to_unsigned(integer(my_cos(3588)),16);
when x"e05" => lut_sig <= to_unsigned(integer(my_cos(3589)),16);
when x"e06" => lut_sig <= to_unsigned(integer(my_cos(3590)),16);
when x"e07" => lut_sig <= to_unsigned(integer(my_cos(3591)),16);
when x"e08" => lut_sig <= to_unsigned(integer(my_cos(3592)),16);
when x"e09" => lut_sig <= to_unsigned(integer(my_cos(3593)),16);
when x"e0a" => lut_sig <= to_unsigned(integer(my_cos(3594)),16);
when x"e0b" => lut_sig <= to_unsigned(integer(my_cos(3595)),16);
when x"e0c" => lut_sig <= to_unsigned(integer(my_cos(3596)),16);
when x"e0d" => lut_sig <= to_unsigned(integer(my_cos(3597)),16);
when x"e0e" => lut_sig <= to_unsigned(integer(my_cos(3598)),16);
when x"e0f" => lut_sig <= to_unsigned(integer(my_cos(3599)),16);
when x"e10" => lut_sig <= to_unsigned(integer(my_cos(3600)),16);
when x"e11" => lut_sig <= to_unsigned(integer(my_cos(3601)),16);
when x"e12" => lut_sig <= to_unsigned(integer(my_cos(3602)),16);
when x"e13" => lut_sig <= to_unsigned(integer(my_cos(3603)),16);
when x"e14" => lut_sig <= to_unsigned(integer(my_cos(3604)),16);
when x"e15" => lut_sig <= to_unsigned(integer(my_cos(3605)),16);
when x"e16" => lut_sig <= to_unsigned(integer(my_cos(3606)),16);
when x"e17" => lut_sig <= to_unsigned(integer(my_cos(3607)),16);
when x"e18" => lut_sig <= to_unsigned(integer(my_cos(3608)),16);
when x"e19" => lut_sig <= to_unsigned(integer(my_cos(3609)),16);
when x"e1a" => lut_sig <= to_unsigned(integer(my_cos(3610)),16);
when x"e1b" => lut_sig <= to_unsigned(integer(my_cos(3611)),16);
when x"e1c" => lut_sig <= to_unsigned(integer(my_cos(3612)),16);
when x"e1d" => lut_sig <= to_unsigned(integer(my_cos(3613)),16);
when x"e1e" => lut_sig <= to_unsigned(integer(my_cos(3614)),16);
when x"e1f" => lut_sig <= to_unsigned(integer(my_cos(3615)),16);
when x"e20" => lut_sig <= to_unsigned(integer(my_cos(3616)),16);
when x"e21" => lut_sig <= to_unsigned(integer(my_cos(3617)),16);
when x"e22" => lut_sig <= to_unsigned(integer(my_cos(3618)),16);
when x"e23" => lut_sig <= to_unsigned(integer(my_cos(3619)),16);
when x"e24" => lut_sig <= to_unsigned(integer(my_cos(3620)),16);
when x"e25" => lut_sig <= to_unsigned(integer(my_cos(3621)),16);
when x"e26" => lut_sig <= to_unsigned(integer(my_cos(3622)),16);
when x"e27" => lut_sig <= to_unsigned(integer(my_cos(3623)),16);
when x"e28" => lut_sig <= to_unsigned(integer(my_cos(3624)),16);
when x"e29" => lut_sig <= to_unsigned(integer(my_cos(3625)),16);
when x"e2a" => lut_sig <= to_unsigned(integer(my_cos(3626)),16);
when x"e2b" => lut_sig <= to_unsigned(integer(my_cos(3627)),16);
when x"e2c" => lut_sig <= to_unsigned(integer(my_cos(3628)),16);
when x"e2d" => lut_sig <= to_unsigned(integer(my_cos(3629)),16);
when x"e2e" => lut_sig <= to_unsigned(integer(my_cos(3630)),16);
when x"e2f" => lut_sig <= to_unsigned(integer(my_cos(3631)),16);
when x"e30" => lut_sig <= to_unsigned(integer(my_cos(3632)),16);
when x"e31" => lut_sig <= to_unsigned(integer(my_cos(3633)),16);
when x"e32" => lut_sig <= to_unsigned(integer(my_cos(3634)),16);
when x"e33" => lut_sig <= to_unsigned(integer(my_cos(3635)),16);
when x"e34" => lut_sig <= to_unsigned(integer(my_cos(3636)),16);
when x"e35" => lut_sig <= to_unsigned(integer(my_cos(3637)),16);
when x"e36" => lut_sig <= to_unsigned(integer(my_cos(3638)),16);
when x"e37" => lut_sig <= to_unsigned(integer(my_cos(3639)),16);
when x"e38" => lut_sig <= to_unsigned(integer(my_cos(3640)),16);
when x"e39" => lut_sig <= to_unsigned(integer(my_cos(3641)),16);
when x"e3a" => lut_sig <= to_unsigned(integer(my_cos(3642)),16);
when x"e3b" => lut_sig <= to_unsigned(integer(my_cos(3643)),16);
when x"e3c" => lut_sig <= to_unsigned(integer(my_cos(3644)),16);
when x"e3d" => lut_sig <= to_unsigned(integer(my_cos(3645)),16);
when x"e3e" => lut_sig <= to_unsigned(integer(my_cos(3646)),16);
when x"e3f" => lut_sig <= to_unsigned(integer(my_cos(3647)),16);
when x"e40" => lut_sig <= to_unsigned(integer(my_cos(3648)),16);
when x"e41" => lut_sig <= to_unsigned(integer(my_cos(3649)),16);
when x"e42" => lut_sig <= to_unsigned(integer(my_cos(3650)),16);
when x"e43" => lut_sig <= to_unsigned(integer(my_cos(3651)),16);
when x"e44" => lut_sig <= to_unsigned(integer(my_cos(3652)),16);
when x"e45" => lut_sig <= to_unsigned(integer(my_cos(3653)),16);
when x"e46" => lut_sig <= to_unsigned(integer(my_cos(3654)),16);
when x"e47" => lut_sig <= to_unsigned(integer(my_cos(3655)),16);
when x"e48" => lut_sig <= to_unsigned(integer(my_cos(3656)),16);
when x"e49" => lut_sig <= to_unsigned(integer(my_cos(3657)),16);
when x"e4a" => lut_sig <= to_unsigned(integer(my_cos(3658)),16);
when x"e4b" => lut_sig <= to_unsigned(integer(my_cos(3659)),16);
when x"e4c" => lut_sig <= to_unsigned(integer(my_cos(3660)),16);
when x"e4d" => lut_sig <= to_unsigned(integer(my_cos(3661)),16);
when x"e4e" => lut_sig <= to_unsigned(integer(my_cos(3662)),16);
when x"e4f" => lut_sig <= to_unsigned(integer(my_cos(3663)),16);
when x"e50" => lut_sig <= to_unsigned(integer(my_cos(3664)),16);
when x"e51" => lut_sig <= to_unsigned(integer(my_cos(3665)),16);
when x"e52" => lut_sig <= to_unsigned(integer(my_cos(3666)),16);
when x"e53" => lut_sig <= to_unsigned(integer(my_cos(3667)),16);
when x"e54" => lut_sig <= to_unsigned(integer(my_cos(3668)),16);
when x"e55" => lut_sig <= to_unsigned(integer(my_cos(3669)),16);
when x"e56" => lut_sig <= to_unsigned(integer(my_cos(3670)),16);
when x"e57" => lut_sig <= to_unsigned(integer(my_cos(3671)),16);
when x"e58" => lut_sig <= to_unsigned(integer(my_cos(3672)),16);
when x"e59" => lut_sig <= to_unsigned(integer(my_cos(3673)),16);
when x"e5a" => lut_sig <= to_unsigned(integer(my_cos(3674)),16);
when x"e5b" => lut_sig <= to_unsigned(integer(my_cos(3675)),16);
when x"e5c" => lut_sig <= to_unsigned(integer(my_cos(3676)),16);
when x"e5d" => lut_sig <= to_unsigned(integer(my_cos(3677)),16);
when x"e5e" => lut_sig <= to_unsigned(integer(my_cos(3678)),16);
when x"e5f" => lut_sig <= to_unsigned(integer(my_cos(3679)),16);
when x"e60" => lut_sig <= to_unsigned(integer(my_cos(3680)),16);
when x"e61" => lut_sig <= to_unsigned(integer(my_cos(3681)),16);
when x"e62" => lut_sig <= to_unsigned(integer(my_cos(3682)),16);
when x"e63" => lut_sig <= to_unsigned(integer(my_cos(3683)),16);
when x"e64" => lut_sig <= to_unsigned(integer(my_cos(3684)),16);
when x"e65" => lut_sig <= to_unsigned(integer(my_cos(3685)),16);
when x"e66" => lut_sig <= to_unsigned(integer(my_cos(3686)),16);
when x"e67" => lut_sig <= to_unsigned(integer(my_cos(3687)),16);
when x"e68" => lut_sig <= to_unsigned(integer(my_cos(3688)),16);
when x"e69" => lut_sig <= to_unsigned(integer(my_cos(3689)),16);
when x"e6a" => lut_sig <= to_unsigned(integer(my_cos(3690)),16);
when x"e6b" => lut_sig <= to_unsigned(integer(my_cos(3691)),16);
when x"e6c" => lut_sig <= to_unsigned(integer(my_cos(3692)),16);
when x"e6d" => lut_sig <= to_unsigned(integer(my_cos(3693)),16);
when x"e6e" => lut_sig <= to_unsigned(integer(my_cos(3694)),16);
when x"e6f" => lut_sig <= to_unsigned(integer(my_cos(3695)),16);
when x"e70" => lut_sig <= to_unsigned(integer(my_cos(3696)),16);
when x"e71" => lut_sig <= to_unsigned(integer(my_cos(3697)),16);
when x"e72" => lut_sig <= to_unsigned(integer(my_cos(3698)),16);
when x"e73" => lut_sig <= to_unsigned(integer(my_cos(3699)),16);
when x"e74" => lut_sig <= to_unsigned(integer(my_cos(3700)),16);
when x"e75" => lut_sig <= to_unsigned(integer(my_cos(3701)),16);
when x"e76" => lut_sig <= to_unsigned(integer(my_cos(3702)),16);
when x"e77" => lut_sig <= to_unsigned(integer(my_cos(3703)),16);
when x"e78" => lut_sig <= to_unsigned(integer(my_cos(3704)),16);
when x"e79" => lut_sig <= to_unsigned(integer(my_cos(3705)),16);
when x"e7a" => lut_sig <= to_unsigned(integer(my_cos(3706)),16);
when x"e7b" => lut_sig <= to_unsigned(integer(my_cos(3707)),16);
when x"e7c" => lut_sig <= to_unsigned(integer(my_cos(3708)),16);
when x"e7d" => lut_sig <= to_unsigned(integer(my_cos(3709)),16);
when x"e7e" => lut_sig <= to_unsigned(integer(my_cos(3710)),16);
when x"e7f" => lut_sig <= to_unsigned(integer(my_cos(3711)),16);
when x"e80" => lut_sig <= to_unsigned(integer(my_cos(3712)),16);
when x"e81" => lut_sig <= to_unsigned(integer(my_cos(3713)),16);
when x"e82" => lut_sig <= to_unsigned(integer(my_cos(3714)),16);
when x"e83" => lut_sig <= to_unsigned(integer(my_cos(3715)),16);
when x"e84" => lut_sig <= to_unsigned(integer(my_cos(3716)),16);
when x"e85" => lut_sig <= to_unsigned(integer(my_cos(3717)),16);
when x"e86" => lut_sig <= to_unsigned(integer(my_cos(3718)),16);
when x"e87" => lut_sig <= to_unsigned(integer(my_cos(3719)),16);
when x"e88" => lut_sig <= to_unsigned(integer(my_cos(3720)),16);
when x"e89" => lut_sig <= to_unsigned(integer(my_cos(3721)),16);
when x"e8a" => lut_sig <= to_unsigned(integer(my_cos(3722)),16);
when x"e8b" => lut_sig <= to_unsigned(integer(my_cos(3723)),16);
when x"e8c" => lut_sig <= to_unsigned(integer(my_cos(3724)),16);
when x"e8d" => lut_sig <= to_unsigned(integer(my_cos(3725)),16);
when x"e8e" => lut_sig <= to_unsigned(integer(my_cos(3726)),16);
when x"e8f" => lut_sig <= to_unsigned(integer(my_cos(3727)),16);
when x"e90" => lut_sig <= to_unsigned(integer(my_cos(3728)),16);
when x"e91" => lut_sig <= to_unsigned(integer(my_cos(3729)),16);
when x"e92" => lut_sig <= to_unsigned(integer(my_cos(3730)),16);
when x"e93" => lut_sig <= to_unsigned(integer(my_cos(3731)),16);
when x"e94" => lut_sig <= to_unsigned(integer(my_cos(3732)),16);
when x"e95" => lut_sig <= to_unsigned(integer(my_cos(3733)),16);
when x"e96" => lut_sig <= to_unsigned(integer(my_cos(3734)),16);
when x"e97" => lut_sig <= to_unsigned(integer(my_cos(3735)),16);
when x"e98" => lut_sig <= to_unsigned(integer(my_cos(3736)),16);
when x"e99" => lut_sig <= to_unsigned(integer(my_cos(3737)),16);
when x"e9a" => lut_sig <= to_unsigned(integer(my_cos(3738)),16);
when x"e9b" => lut_sig <= to_unsigned(integer(my_cos(3739)),16);
when x"e9c" => lut_sig <= to_unsigned(integer(my_cos(3740)),16);
when x"e9d" => lut_sig <= to_unsigned(integer(my_cos(3741)),16);
when x"e9e" => lut_sig <= to_unsigned(integer(my_cos(3742)),16);
when x"e9f" => lut_sig <= to_unsigned(integer(my_cos(3743)),16);
when x"ea0" => lut_sig <= to_unsigned(integer(my_cos(3744)),16);
when x"ea1" => lut_sig <= to_unsigned(integer(my_cos(3745)),16);
when x"ea2" => lut_sig <= to_unsigned(integer(my_cos(3746)),16);
when x"ea3" => lut_sig <= to_unsigned(integer(my_cos(3747)),16);
when x"ea4" => lut_sig <= to_unsigned(integer(my_cos(3748)),16);
when x"ea5" => lut_sig <= to_unsigned(integer(my_cos(3749)),16);
when x"ea6" => lut_sig <= to_unsigned(integer(my_cos(3750)),16);
when x"ea7" => lut_sig <= to_unsigned(integer(my_cos(3751)),16);
when x"ea8" => lut_sig <= to_unsigned(integer(my_cos(3752)),16);
when x"ea9" => lut_sig <= to_unsigned(integer(my_cos(3753)),16);
when x"eaa" => lut_sig <= to_unsigned(integer(my_cos(3754)),16);
when x"eab" => lut_sig <= to_unsigned(integer(my_cos(3755)),16);
when x"eac" => lut_sig <= to_unsigned(integer(my_cos(3756)),16);
when x"ead" => lut_sig <= to_unsigned(integer(my_cos(3757)),16);
when x"eae" => lut_sig <= to_unsigned(integer(my_cos(3758)),16);
when x"eaf" => lut_sig <= to_unsigned(integer(my_cos(3759)),16);
when x"eb0" => lut_sig <= to_unsigned(integer(my_cos(3760)),16);
when x"eb1" => lut_sig <= to_unsigned(integer(my_cos(3761)),16);
when x"eb2" => lut_sig <= to_unsigned(integer(my_cos(3762)),16);
when x"eb3" => lut_sig <= to_unsigned(integer(my_cos(3763)),16);
when x"eb4" => lut_sig <= to_unsigned(integer(my_cos(3764)),16);
when x"eb5" => lut_sig <= to_unsigned(integer(my_cos(3765)),16);
when x"eb6" => lut_sig <= to_unsigned(integer(my_cos(3766)),16);
when x"eb7" => lut_sig <= to_unsigned(integer(my_cos(3767)),16);
when x"eb8" => lut_sig <= to_unsigned(integer(my_cos(3768)),16);
when x"eb9" => lut_sig <= to_unsigned(integer(my_cos(3769)),16);
when x"eba" => lut_sig <= to_unsigned(integer(my_cos(3770)),16);
when x"ebb" => lut_sig <= to_unsigned(integer(my_cos(3771)),16);
when x"ebc" => lut_sig <= to_unsigned(integer(my_cos(3772)),16);
when x"ebd" => lut_sig <= to_unsigned(integer(my_cos(3773)),16);
when x"ebe" => lut_sig <= to_unsigned(integer(my_cos(3774)),16);
when x"ebf" => lut_sig <= to_unsigned(integer(my_cos(3775)),16);
when x"ec0" => lut_sig <= to_unsigned(integer(my_cos(3776)),16);
when x"ec1" => lut_sig <= to_unsigned(integer(my_cos(3777)),16);
when x"ec2" => lut_sig <= to_unsigned(integer(my_cos(3778)),16);
when x"ec3" => lut_sig <= to_unsigned(integer(my_cos(3779)),16);
when x"ec4" => lut_sig <= to_unsigned(integer(my_cos(3780)),16);
when x"ec5" => lut_sig <= to_unsigned(integer(my_cos(3781)),16);
when x"ec6" => lut_sig <= to_unsigned(integer(my_cos(3782)),16);
when x"ec7" => lut_sig <= to_unsigned(integer(my_cos(3783)),16);
when x"ec8" => lut_sig <= to_unsigned(integer(my_cos(3784)),16);
when x"ec9" => lut_sig <= to_unsigned(integer(my_cos(3785)),16);
when x"eca" => lut_sig <= to_unsigned(integer(my_cos(3786)),16);
when x"ecb" => lut_sig <= to_unsigned(integer(my_cos(3787)),16);
when x"ecc" => lut_sig <= to_unsigned(integer(my_cos(3788)),16);
when x"ecd" => lut_sig <= to_unsigned(integer(my_cos(3789)),16);
when x"ece" => lut_sig <= to_unsigned(integer(my_cos(3790)),16);
when x"ecf" => lut_sig <= to_unsigned(integer(my_cos(3791)),16);
when x"ed0" => lut_sig <= to_unsigned(integer(my_cos(3792)),16);
when x"ed1" => lut_sig <= to_unsigned(integer(my_cos(3793)),16);
when x"ed2" => lut_sig <= to_unsigned(integer(my_cos(3794)),16);
when x"ed3" => lut_sig <= to_unsigned(integer(my_cos(3795)),16);
when x"ed4" => lut_sig <= to_unsigned(integer(my_cos(3796)),16);
when x"ed5" => lut_sig <= to_unsigned(integer(my_cos(3797)),16);
when x"ed6" => lut_sig <= to_unsigned(integer(my_cos(3798)),16);
when x"ed7" => lut_sig <= to_unsigned(integer(my_cos(3799)),16);
when x"ed8" => lut_sig <= to_unsigned(integer(my_cos(3800)),16);
when x"ed9" => lut_sig <= to_unsigned(integer(my_cos(3801)),16);
when x"eda" => lut_sig <= to_unsigned(integer(my_cos(3802)),16);
when x"edb" => lut_sig <= to_unsigned(integer(my_cos(3803)),16);
when x"edc" => lut_sig <= to_unsigned(integer(my_cos(3804)),16);
when x"edd" => lut_sig <= to_unsigned(integer(my_cos(3805)),16);
when x"ede" => lut_sig <= to_unsigned(integer(my_cos(3806)),16);
when x"edf" => lut_sig <= to_unsigned(integer(my_cos(3807)),16);
when x"ee0" => lut_sig <= to_unsigned(integer(my_cos(3808)),16);
when x"ee1" => lut_sig <= to_unsigned(integer(my_cos(3809)),16);
when x"ee2" => lut_sig <= to_unsigned(integer(my_cos(3810)),16);
when x"ee3" => lut_sig <= to_unsigned(integer(my_cos(3811)),16);
when x"ee4" => lut_sig <= to_unsigned(integer(my_cos(3812)),16);
when x"ee5" => lut_sig <= to_unsigned(integer(my_cos(3813)),16);
when x"ee6" => lut_sig <= to_unsigned(integer(my_cos(3814)),16);
when x"ee7" => lut_sig <= to_unsigned(integer(my_cos(3815)),16);
when x"ee8" => lut_sig <= to_unsigned(integer(my_cos(3816)),16);
when x"ee9" => lut_sig <= to_unsigned(integer(my_cos(3817)),16);
when x"eea" => lut_sig <= to_unsigned(integer(my_cos(3818)),16);
when x"eeb" => lut_sig <= to_unsigned(integer(my_cos(3819)),16);
when x"eec" => lut_sig <= to_unsigned(integer(my_cos(3820)),16);
when x"eed" => lut_sig <= to_unsigned(integer(my_cos(3821)),16);
when x"eee" => lut_sig <= to_unsigned(integer(my_cos(3822)),16);
when x"eef" => lut_sig <= to_unsigned(integer(my_cos(3823)),16);
when x"ef0" => lut_sig <= to_unsigned(integer(my_cos(3824)),16);
when x"ef1" => lut_sig <= to_unsigned(integer(my_cos(3825)),16);
when x"ef2" => lut_sig <= to_unsigned(integer(my_cos(3826)),16);
when x"ef3" => lut_sig <= to_unsigned(integer(my_cos(3827)),16);
when x"ef4" => lut_sig <= to_unsigned(integer(my_cos(3828)),16);
when x"ef5" => lut_sig <= to_unsigned(integer(my_cos(3829)),16);
when x"ef6" => lut_sig <= to_unsigned(integer(my_cos(3830)),16);
when x"ef7" => lut_sig <= to_unsigned(integer(my_cos(3831)),16);
when x"ef8" => lut_sig <= to_unsigned(integer(my_cos(3832)),16);
when x"ef9" => lut_sig <= to_unsigned(integer(my_cos(3833)),16);
when x"efa" => lut_sig <= to_unsigned(integer(my_cos(3834)),16);
when x"efb" => lut_sig <= to_unsigned(integer(my_cos(3835)),16);
when x"efc" => lut_sig <= to_unsigned(integer(my_cos(3836)),16);
when x"efd" => lut_sig <= to_unsigned(integer(my_cos(3837)),16);
when x"efe" => lut_sig <= to_unsigned(integer(my_cos(3838)),16);
when x"eff" => lut_sig <= to_unsigned(integer(my_cos(3839)),16);
when x"f00" => lut_sig <= to_unsigned(integer(my_cos(3840)),16);
when x"f01" => lut_sig <= to_unsigned(integer(my_cos(3841)),16);
when x"f02" => lut_sig <= to_unsigned(integer(my_cos(3842)),16);
when x"f03" => lut_sig <= to_unsigned(integer(my_cos(3843)),16);
when x"f04" => lut_sig <= to_unsigned(integer(my_cos(3844)),16);
when x"f05" => lut_sig <= to_unsigned(integer(my_cos(3845)),16);
when x"f06" => lut_sig <= to_unsigned(integer(my_cos(3846)),16);
when x"f07" => lut_sig <= to_unsigned(integer(my_cos(3847)),16);
when x"f08" => lut_sig <= to_unsigned(integer(my_cos(3848)),16);
when x"f09" => lut_sig <= to_unsigned(integer(my_cos(3849)),16);
when x"f0a" => lut_sig <= to_unsigned(integer(my_cos(3850)),16);
when x"f0b" => lut_sig <= to_unsigned(integer(my_cos(3851)),16);
when x"f0c" => lut_sig <= to_unsigned(integer(my_cos(3852)),16);
when x"f0d" => lut_sig <= to_unsigned(integer(my_cos(3853)),16);
when x"f0e" => lut_sig <= to_unsigned(integer(my_cos(3854)),16);
when x"f0f" => lut_sig <= to_unsigned(integer(my_cos(3855)),16);
when x"f10" => lut_sig <= to_unsigned(integer(my_cos(3856)),16);
when x"f11" => lut_sig <= to_unsigned(integer(my_cos(3857)),16);
when x"f12" => lut_sig <= to_unsigned(integer(my_cos(3858)),16);
when x"f13" => lut_sig <= to_unsigned(integer(my_cos(3859)),16);
when x"f14" => lut_sig <= to_unsigned(integer(my_cos(3860)),16);
when x"f15" => lut_sig <= to_unsigned(integer(my_cos(3861)),16);
when x"f16" => lut_sig <= to_unsigned(integer(my_cos(3862)),16);
when x"f17" => lut_sig <= to_unsigned(integer(my_cos(3863)),16);
when x"f18" => lut_sig <= to_unsigned(integer(my_cos(3864)),16);
when x"f19" => lut_sig <= to_unsigned(integer(my_cos(3865)),16);
when x"f1a" => lut_sig <= to_unsigned(integer(my_cos(3866)),16);
when x"f1b" => lut_sig <= to_unsigned(integer(my_cos(3867)),16);
when x"f1c" => lut_sig <= to_unsigned(integer(my_cos(3868)),16);
when x"f1d" => lut_sig <= to_unsigned(integer(my_cos(3869)),16);
when x"f1e" => lut_sig <= to_unsigned(integer(my_cos(3870)),16);
when x"f1f" => lut_sig <= to_unsigned(integer(my_cos(3871)),16);
when x"f20" => lut_sig <= to_unsigned(integer(my_cos(3872)),16);
when x"f21" => lut_sig <= to_unsigned(integer(my_cos(3873)),16);
when x"f22" => lut_sig <= to_unsigned(integer(my_cos(3874)),16);
when x"f23" => lut_sig <= to_unsigned(integer(my_cos(3875)),16);
when x"f24" => lut_sig <= to_unsigned(integer(my_cos(3876)),16);
when x"f25" => lut_sig <= to_unsigned(integer(my_cos(3877)),16);
when x"f26" => lut_sig <= to_unsigned(integer(my_cos(3878)),16);
when x"f27" => lut_sig <= to_unsigned(integer(my_cos(3879)),16);
when x"f28" => lut_sig <= to_unsigned(integer(my_cos(3880)),16);
when x"f29" => lut_sig <= to_unsigned(integer(my_cos(3881)),16);
when x"f2a" => lut_sig <= to_unsigned(integer(my_cos(3882)),16);
when x"f2b" => lut_sig <= to_unsigned(integer(my_cos(3883)),16);
when x"f2c" => lut_sig <= to_unsigned(integer(my_cos(3884)),16);
when x"f2d" => lut_sig <= to_unsigned(integer(my_cos(3885)),16);
when x"f2e" => lut_sig <= to_unsigned(integer(my_cos(3886)),16);
when x"f2f" => lut_sig <= to_unsigned(integer(my_cos(3887)),16);
when x"f30" => lut_sig <= to_unsigned(integer(my_cos(3888)),16);
when x"f31" => lut_sig <= to_unsigned(integer(my_cos(3889)),16);
when x"f32" => lut_sig <= to_unsigned(integer(my_cos(3890)),16);
when x"f33" => lut_sig <= to_unsigned(integer(my_cos(3891)),16);
when x"f34" => lut_sig <= to_unsigned(integer(my_cos(3892)),16);
when x"f35" => lut_sig <= to_unsigned(integer(my_cos(3893)),16);
when x"f36" => lut_sig <= to_unsigned(integer(my_cos(3894)),16);
when x"f37" => lut_sig <= to_unsigned(integer(my_cos(3895)),16);
when x"f38" => lut_sig <= to_unsigned(integer(my_cos(3896)),16);
when x"f39" => lut_sig <= to_unsigned(integer(my_cos(3897)),16);
when x"f3a" => lut_sig <= to_unsigned(integer(my_cos(3898)),16);
when x"f3b" => lut_sig <= to_unsigned(integer(my_cos(3899)),16);
when x"f3c" => lut_sig <= to_unsigned(integer(my_cos(3900)),16);
when x"f3d" => lut_sig <= to_unsigned(integer(my_cos(3901)),16);
when x"f3e" => lut_sig <= to_unsigned(integer(my_cos(3902)),16);
when x"f3f" => lut_sig <= to_unsigned(integer(my_cos(3903)),16);
when x"f40" => lut_sig <= to_unsigned(integer(my_cos(3904)),16);
when x"f41" => lut_sig <= to_unsigned(integer(my_cos(3905)),16);
when x"f42" => lut_sig <= to_unsigned(integer(my_cos(3906)),16);
when x"f43" => lut_sig <= to_unsigned(integer(my_cos(3907)),16);
when x"f44" => lut_sig <= to_unsigned(integer(my_cos(3908)),16);
when x"f45" => lut_sig <= to_unsigned(integer(my_cos(3909)),16);
when x"f46" => lut_sig <= to_unsigned(integer(my_cos(3910)),16);
when x"f47" => lut_sig <= to_unsigned(integer(my_cos(3911)),16);
when x"f48" => lut_sig <= to_unsigned(integer(my_cos(3912)),16);
when x"f49" => lut_sig <= to_unsigned(integer(my_cos(3913)),16);
when x"f4a" => lut_sig <= to_unsigned(integer(my_cos(3914)),16);
when x"f4b" => lut_sig <= to_unsigned(integer(my_cos(3915)),16);
when x"f4c" => lut_sig <= to_unsigned(integer(my_cos(3916)),16);
when x"f4d" => lut_sig <= to_unsigned(integer(my_cos(3917)),16);
when x"f4e" => lut_sig <= to_unsigned(integer(my_cos(3918)),16);
when x"f4f" => lut_sig <= to_unsigned(integer(my_cos(3919)),16);
when x"f50" => lut_sig <= to_unsigned(integer(my_cos(3920)),16);
when x"f51" => lut_sig <= to_unsigned(integer(my_cos(3921)),16);
when x"f52" => lut_sig <= to_unsigned(integer(my_cos(3922)),16);
when x"f53" => lut_sig <= to_unsigned(integer(my_cos(3923)),16);
when x"f54" => lut_sig <= to_unsigned(integer(my_cos(3924)),16);
when x"f55" => lut_sig <= to_unsigned(integer(my_cos(3925)),16);
when x"f56" => lut_sig <= to_unsigned(integer(my_cos(3926)),16);
when x"f57" => lut_sig <= to_unsigned(integer(my_cos(3927)),16);
when x"f58" => lut_sig <= to_unsigned(integer(my_cos(3928)),16);
when x"f59" => lut_sig <= to_unsigned(integer(my_cos(3929)),16);
when x"f5a" => lut_sig <= to_unsigned(integer(my_cos(3930)),16);
when x"f5b" => lut_sig <= to_unsigned(integer(my_cos(3931)),16);
when x"f5c" => lut_sig <= to_unsigned(integer(my_cos(3932)),16);
when x"f5d" => lut_sig <= to_unsigned(integer(my_cos(3933)),16);
when x"f5e" => lut_sig <= to_unsigned(integer(my_cos(3934)),16);
when x"f5f" => lut_sig <= to_unsigned(integer(my_cos(3935)),16);
when x"f60" => lut_sig <= to_unsigned(integer(my_cos(3936)),16);
when x"f61" => lut_sig <= to_unsigned(integer(my_cos(3937)),16);
when x"f62" => lut_sig <= to_unsigned(integer(my_cos(3938)),16);
when x"f63" => lut_sig <= to_unsigned(integer(my_cos(3939)),16);
when x"f64" => lut_sig <= to_unsigned(integer(my_cos(3940)),16);
when x"f65" => lut_sig <= to_unsigned(integer(my_cos(3941)),16);
when x"f66" => lut_sig <= to_unsigned(integer(my_cos(3942)),16);
when x"f67" => lut_sig <= to_unsigned(integer(my_cos(3943)),16);
when x"f68" => lut_sig <= to_unsigned(integer(my_cos(3944)),16);
when x"f69" => lut_sig <= to_unsigned(integer(my_cos(3945)),16);
when x"f6a" => lut_sig <= to_unsigned(integer(my_cos(3946)),16);
when x"f6b" => lut_sig <= to_unsigned(integer(my_cos(3947)),16);
when x"f6c" => lut_sig <= to_unsigned(integer(my_cos(3948)),16);
when x"f6d" => lut_sig <= to_unsigned(integer(my_cos(3949)),16);
when x"f6e" => lut_sig <= to_unsigned(integer(my_cos(3950)),16);
when x"f6f" => lut_sig <= to_unsigned(integer(my_cos(3951)),16);
when x"f70" => lut_sig <= to_unsigned(integer(my_cos(3952)),16);
when x"f71" => lut_sig <= to_unsigned(integer(my_cos(3953)),16);
when x"f72" => lut_sig <= to_unsigned(integer(my_cos(3954)),16);
when x"f73" => lut_sig <= to_unsigned(integer(my_cos(3955)),16);
when x"f74" => lut_sig <= to_unsigned(integer(my_cos(3956)),16);
when x"f75" => lut_sig <= to_unsigned(integer(my_cos(3957)),16);
when x"f76" => lut_sig <= to_unsigned(integer(my_cos(3958)),16);
when x"f77" => lut_sig <= to_unsigned(integer(my_cos(3959)),16);
when x"f78" => lut_sig <= to_unsigned(integer(my_cos(3960)),16);
when x"f79" => lut_sig <= to_unsigned(integer(my_cos(3961)),16);
when x"f7a" => lut_sig <= to_unsigned(integer(my_cos(3962)),16);
when x"f7b" => lut_sig <= to_unsigned(integer(my_cos(3963)),16);
when x"f7c" => lut_sig <= to_unsigned(integer(my_cos(3964)),16);
when x"f7d" => lut_sig <= to_unsigned(integer(my_cos(3965)),16);
when x"f7e" => lut_sig <= to_unsigned(integer(my_cos(3966)),16);
when x"f7f" => lut_sig <= to_unsigned(integer(my_cos(3967)),16);
when x"f80" => lut_sig <= to_unsigned(integer(my_cos(3968)),16);
when x"f81" => lut_sig <= to_unsigned(integer(my_cos(3969)),16);
when x"f82" => lut_sig <= to_unsigned(integer(my_cos(3970)),16);
when x"f83" => lut_sig <= to_unsigned(integer(my_cos(3971)),16);
when x"f84" => lut_sig <= to_unsigned(integer(my_cos(3972)),16);
when x"f85" => lut_sig <= to_unsigned(integer(my_cos(3973)),16);
when x"f86" => lut_sig <= to_unsigned(integer(my_cos(3974)),16);
when x"f87" => lut_sig <= to_unsigned(integer(my_cos(3975)),16);
when x"f88" => lut_sig <= to_unsigned(integer(my_cos(3976)),16);
when x"f89" => lut_sig <= to_unsigned(integer(my_cos(3977)),16);
when x"f8a" => lut_sig <= to_unsigned(integer(my_cos(3978)),16);
when x"f8b" => lut_sig <= to_unsigned(integer(my_cos(3979)),16);
when x"f8c" => lut_sig <= to_unsigned(integer(my_cos(3980)),16);
when x"f8d" => lut_sig <= to_unsigned(integer(my_cos(3981)),16);
when x"f8e" => lut_sig <= to_unsigned(integer(my_cos(3982)),16);
when x"f8f" => lut_sig <= to_unsigned(integer(my_cos(3983)),16);
when x"f90" => lut_sig <= to_unsigned(integer(my_cos(3984)),16);
when x"f91" => lut_sig <= to_unsigned(integer(my_cos(3985)),16);
when x"f92" => lut_sig <= to_unsigned(integer(my_cos(3986)),16);
when x"f93" => lut_sig <= to_unsigned(integer(my_cos(3987)),16);
when x"f94" => lut_sig <= to_unsigned(integer(my_cos(3988)),16);
when x"f95" => lut_sig <= to_unsigned(integer(my_cos(3989)),16);
when x"f96" => lut_sig <= to_unsigned(integer(my_cos(3990)),16);
when x"f97" => lut_sig <= to_unsigned(integer(my_cos(3991)),16);
when x"f98" => lut_sig <= to_unsigned(integer(my_cos(3992)),16);
when x"f99" => lut_sig <= to_unsigned(integer(my_cos(3993)),16);
when x"f9a" => lut_sig <= to_unsigned(integer(my_cos(3994)),16);
when x"f9b" => lut_sig <= to_unsigned(integer(my_cos(3995)),16);
when x"f9c" => lut_sig <= to_unsigned(integer(my_cos(3996)),16);
when x"f9d" => lut_sig <= to_unsigned(integer(my_cos(3997)),16);
when x"f9e" => lut_sig <= to_unsigned(integer(my_cos(3998)),16);
when x"f9f" => lut_sig <= to_unsigned(integer(my_cos(3999)),16);
when x"fa0" => lut_sig <= to_unsigned(integer(my_cos(4000)),16);
when x"fa1" => lut_sig <= to_unsigned(integer(my_cos(4001)),16);
when x"fa2" => lut_sig <= to_unsigned(integer(my_cos(4002)),16);
when x"fa3" => lut_sig <= to_unsigned(integer(my_cos(4003)),16);
when x"fa4" => lut_sig <= to_unsigned(integer(my_cos(4004)),16);
when x"fa5" => lut_sig <= to_unsigned(integer(my_cos(4005)),16);
when x"fa6" => lut_sig <= to_unsigned(integer(my_cos(4006)),16);
when x"fa7" => lut_sig <= to_unsigned(integer(my_cos(4007)),16);
when x"fa8" => lut_sig <= to_unsigned(integer(my_cos(4008)),16);
when x"fa9" => lut_sig <= to_unsigned(integer(my_cos(4009)),16);
when x"faa" => lut_sig <= to_unsigned(integer(my_cos(4010)),16);
when x"fab" => lut_sig <= to_unsigned(integer(my_cos(4011)),16);
when x"fac" => lut_sig <= to_unsigned(integer(my_cos(4012)),16);
when x"fad" => lut_sig <= to_unsigned(integer(my_cos(4013)),16);
when x"fae" => lut_sig <= to_unsigned(integer(my_cos(4014)),16);
when x"faf" => lut_sig <= to_unsigned(integer(my_cos(4015)),16);
when x"fb0" => lut_sig <= to_unsigned(integer(my_cos(4016)),16);
when x"fb1" => lut_sig <= to_unsigned(integer(my_cos(4017)),16);
when x"fb2" => lut_sig <= to_unsigned(integer(my_cos(4018)),16);
when x"fb3" => lut_sig <= to_unsigned(integer(my_cos(4019)),16);
when x"fb4" => lut_sig <= to_unsigned(integer(my_cos(4020)),16);
when x"fb5" => lut_sig <= to_unsigned(integer(my_cos(4021)),16);
when x"fb6" => lut_sig <= to_unsigned(integer(my_cos(4022)),16);
when x"fb7" => lut_sig <= to_unsigned(integer(my_cos(4023)),16);
when x"fb8" => lut_sig <= to_unsigned(integer(my_cos(4024)),16);
when x"fb9" => lut_sig <= to_unsigned(integer(my_cos(4025)),16);
when x"fba" => lut_sig <= to_unsigned(integer(my_cos(4026)),16);
when x"fbb" => lut_sig <= to_unsigned(integer(my_cos(4027)),16);
when x"fbc" => lut_sig <= to_unsigned(integer(my_cos(4028)),16);
when x"fbd" => lut_sig <= to_unsigned(integer(my_cos(4029)),16);
when x"fbe" => lut_sig <= to_unsigned(integer(my_cos(4030)),16);
when x"fbf" => lut_sig <= to_unsigned(integer(my_cos(4031)),16);
when x"fc0" => lut_sig <= to_unsigned(integer(my_cos(4032)),16);
when x"fc1" => lut_sig <= to_unsigned(integer(my_cos(4033)),16);
when x"fc2" => lut_sig <= to_unsigned(integer(my_cos(4034)),16);
when x"fc3" => lut_sig <= to_unsigned(integer(my_cos(4035)),16);
when x"fc4" => lut_sig <= to_unsigned(integer(my_cos(4036)),16);
when x"fc5" => lut_sig <= to_unsigned(integer(my_cos(4037)),16);
when x"fc6" => lut_sig <= to_unsigned(integer(my_cos(4038)),16);
when x"fc7" => lut_sig <= to_unsigned(integer(my_cos(4039)),16);
when x"fc8" => lut_sig <= to_unsigned(integer(my_cos(4040)),16);
when x"fc9" => lut_sig <= to_unsigned(integer(my_cos(4041)),16);
when x"fca" => lut_sig <= to_unsigned(integer(my_cos(4042)),16);
when x"fcb" => lut_sig <= to_unsigned(integer(my_cos(4043)),16);
when x"fcc" => lut_sig <= to_unsigned(integer(my_cos(4044)),16);
when x"fcd" => lut_sig <= to_unsigned(integer(my_cos(4045)),16);
when x"fce" => lut_sig <= to_unsigned(integer(my_cos(4046)),16);
when x"fcf" => lut_sig <= to_unsigned(integer(my_cos(4047)),16);
when x"fd0" => lut_sig <= to_unsigned(integer(my_cos(4048)),16);
when x"fd1" => lut_sig <= to_unsigned(integer(my_cos(4049)),16);
when x"fd2" => lut_sig <= to_unsigned(integer(my_cos(4050)),16);
when x"fd3" => lut_sig <= to_unsigned(integer(my_cos(4051)),16);
when x"fd4" => lut_sig <= to_unsigned(integer(my_cos(4052)),16);
when x"fd5" => lut_sig <= to_unsigned(integer(my_cos(4053)),16);
when x"fd6" => lut_sig <= to_unsigned(integer(my_cos(4054)),16);
when x"fd7" => lut_sig <= to_unsigned(integer(my_cos(4055)),16);
when x"fd8" => lut_sig <= to_unsigned(integer(my_cos(4056)),16);
when x"fd9" => lut_sig <= to_unsigned(integer(my_cos(4057)),16);
when x"fda" => lut_sig <= to_unsigned(integer(my_cos(4058)),16);
when x"fdb" => lut_sig <= to_unsigned(integer(my_cos(4059)),16);
when x"fdc" => lut_sig <= to_unsigned(integer(my_cos(4060)),16);
when x"fdd" => lut_sig <= to_unsigned(integer(my_cos(4061)),16);
when x"fde" => lut_sig <= to_unsigned(integer(my_cos(4062)),16);
when x"fdf" => lut_sig <= to_unsigned(integer(my_cos(4063)),16);
when x"fe0" => lut_sig <= to_unsigned(integer(my_cos(4064)),16);
when x"fe1" => lut_sig <= to_unsigned(integer(my_cos(4065)),16);
when x"fe2" => lut_sig <= to_unsigned(integer(my_cos(4066)),16);
when x"fe3" => lut_sig <= to_unsigned(integer(my_cos(4067)),16);
when x"fe4" => lut_sig <= to_unsigned(integer(my_cos(4068)),16);
when x"fe5" => lut_sig <= to_unsigned(integer(my_cos(4069)),16);
when x"fe6" => lut_sig <= to_unsigned(integer(my_cos(4070)),16);
when x"fe7" => lut_sig <= to_unsigned(integer(my_cos(4071)),16);
when x"fe8" => lut_sig <= to_unsigned(integer(my_cos(4072)),16);
when x"fe9" => lut_sig <= to_unsigned(integer(my_cos(4073)),16);
when x"fea" => lut_sig <= to_unsigned(integer(my_cos(4074)),16);
when x"feb" => lut_sig <= to_unsigned(integer(my_cos(4075)),16);
when x"fec" => lut_sig <= to_unsigned(integer(my_cos(4076)),16);
when x"fed" => lut_sig <= to_unsigned(integer(my_cos(4077)),16);
when x"fee" => lut_sig <= to_unsigned(integer(my_cos(4078)),16);
when x"fef" => lut_sig <= to_unsigned(integer(my_cos(4079)),16);
when x"ff0" => lut_sig <= to_unsigned(integer(my_cos(4080)),16);
when x"ff1" => lut_sig <= to_unsigned(integer(my_cos(4081)),16);
when x"ff2" => lut_sig <= to_unsigned(integer(my_cos(4082)),16);
when x"ff3" => lut_sig <= to_unsigned(integer(my_cos(4083)),16);
when x"ff4" => lut_sig <= to_unsigned(integer(my_cos(4084)),16);
when x"ff5" => lut_sig <= to_unsigned(integer(my_cos(4085)),16);
when x"ff6" => lut_sig <= to_unsigned(integer(my_cos(4086)),16);
when x"ff7" => lut_sig <= to_unsigned(integer(my_cos(4087)),16);
when x"ff8" => lut_sig <= to_unsigned(integer(my_cos(4088)),16);
when x"ff9" => lut_sig <= to_unsigned(integer(my_cos(4089)),16);
when x"ffa" => lut_sig <= to_unsigned(integer(my_cos(4090)),16);
when x"ffb" => lut_sig <= to_unsigned(integer(my_cos(4091)),16);
when x"ffc" => lut_sig <= to_unsigned(integer(my_cos(4092)),16);
when x"ffd" => lut_sig <= to_unsigned(integer(my_cos(4093)),16);
when x"ffe" => lut_sig <= to_unsigned(integer(my_cos(4094)),16);
when x"fff" => lut_sig <= to_unsigned(integer(my_cos(4095)),16);
                    when others => lut_sig <= "0000000000000000";
                end case;
            end process;
end Behavioral;
