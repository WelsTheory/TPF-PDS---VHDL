library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity sine_lut_prueba is
    Port (
        clk: in STD_LOGIC;
        rst: in STD_LOGIC;
        sine: out STD_LOGIC_VECTOR(15 downto 0)
    );
end entity;

architecture Behavioral of sine_lut_prueba is
    
    type mem is array(0 to 99) of real;
    constant my_rom: mem := (
        0=>750.0,
1=>797.5679397424234,
2=>844.944340180312,
3=>891.9384332703077,
4=>938.3609903858094,
5=>984.0250842738653,
6=>1028.7468417452455,
7=>1072.3461840668788,
8=>1114.6475520753515,
9=>1155.4806130916982,
10=>1194.6809467909804,
11=>1232.0907072649045,
12=>1267.559258611584,
13=>1300.94378149315,
14=>1332.1098482188177,
15=>1360.9319640377516,
16=>1387.2940724621358,
17=>1411.0900225856867,
18=>1432.2239965158888,
19=>1450.61089519883,
20=>1466.1766810830554,
21=>1478.8586762426562,
22=>1488.6058147591561,
23=>1495.3788483459407,
24=>1499.150504387256,
25=>1499.9055957554065,
26=>1497.6410819639568,
27=>1492.3660814106995,
28=>1484.101834661084,
29=>1472.8816189199565,
30=>1458.7506140360015,
31=>1441.765720578436,
32=>1421.995330718502,
33=>1399.519052838329,
34=>1374.4273909760784,
35=>1346.821380398124,
36=>1316.8121807656937,
37=>1284.520628534147,
38=>1250.076750387219,
39=>1213.6192396654537,
40=>1175.2948978970778,
41=>1135.2580436800547,
42=>1093.6698912955578,
43=>1050.6979015549603,
44=>1006.5151074942514,
45=>961.2994176310723,
46=>915.2328995899053,
47=>868.5010469800121,
48=>821.2920324781371,
49=>773.7959501235507,
50=>726.2040498764491,
51=>678.7079675218627,
52=>631.4989530199874,
53=>584.7671004100946,
54=>538.7005823689276,
55=>493.4848925057485,
56=>449.30209844503935,
57=>406.330108704442,
58=>364.7419563199454,
59=>324.7051021029218,
60=>286.38076033454604,
61=>249.9232496127811,
62=>215.47937146585275,
63=>183.18781923430595,
64=>153.17861960187588,
65=>125.57260902392159,
66=>100.48094716167088,
67=>78.00466928149797,
68=>58.23427942156377,
69=>41.24938596399875,
70=>27.118381080043378,
71=>15.898165338915987,
72=>7.633918589300492,
73=>2.3589180360431783,
74=>0.09440424459364749,
75=>0.8494956127440219,
76=>4.6211516540594175,
77=>11.394185240843854,
78=>21.141323757343798,
79=>33.82331891694457,
80=>49.38910480117022,
81=>67.77600348411136,
82=>88.90997741431352,
83=>112.70592753786423,
84=>139.06803596224813,
85=>167.89015178118257,
86=>199.0562185068501,
87=>232.44074138841643,
88=>267.9092927350958,
89=>305.31905320901984,
90=>344.5193869083019,
91=>385.3524479246484,
92=>427.6538159331216,
93=>471.25315825475457,
94=>515.9749157261354,
95=>561.6390096141904,
96=>608.061566729692,
97=>655.0556598196882,
98=>702.4320602575766,
99=>749.9999999999998
    );

signal lut_sig : unsigned(15 downto 0);
signal state : STD_LOGIC;
begin 

sine <= STD_LOGIC_VECTOR(lut_sig);-- when state = '0' else
        --STD_LOGIC_VECTOR(2-lut_sig);
process(clk,rst) is
variable cnt : integer range 0 to 100;
begin
    if rst = '0' then
        cnt := 0;
        state <= '0'; 
        lut_sig <= (others=>'0');
    elsif rising_edge(clk) then
        lut_sig <= to_unsigned(integer(my_rom(cnt)),16);
        if cnt > 98 then
            cnt := 0;
            state <= not state;
        else
            cnt := cnt + 1;
        end if;
    end if;
end process;

end Behavioral;
